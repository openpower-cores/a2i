library ieee;
use ieee.std_logic_1164.all;

package vcomponents is
  component BRAM_TDP_MACRO
    generic (
      BRAM_SIZE           : string;
      DEVICE              : string;
      DOA_REG             : integer;
      DOB_REG             : integer;
      INIT_A              : bit_vector;
      INIT_B              : bit_vector;
      INIT_FILE           : string;
      READ_WIDTH_A        : integer;
      READ_WIDTH_B        : integer;
      SIM_COLLISION_CHECK : string;
      SRVAL_A             : bit_vector;
      SRVAL_B             : bit_vector;
      WRITE_MODE_A        : string;
      WRITE_MODE_B        : string;
      WRITE_WIDTH_A       : integer;
      WRITE_WIDTH_B       : integer;
      INIT_00             : bit_vector;
      INIT_01             : bit_vector;
      INIT_02             : bit_vector;
      INIT_03             : bit_vector;
      INIT_04             : bit_vector;
      INIT_05             : bit_vector;
      INIT_06             : bit_vector;
      INIT_07             : bit_vector;
      INIT_08             : bit_vector;
      INIT_09             : bit_vector;
      INIT_0A             : bit_vector;
      INIT_0B             : bit_vector;
      INIT_0C             : bit_vector;
      INIT_0D             : bit_vector;
      INIT_0E             : bit_vector;
      INIT_0F             : bit_vector;
      INIT_10             : bit_vector;
      INIT_11             : bit_vector;
      INIT_12             : bit_vector;
      INIT_13             : bit_vector;
      INIT_14             : bit_vector;
      INIT_15             : bit_vector;
      INIT_16             : bit_vector;
      INIT_17             : bit_vector;
      INIT_18             : bit_vector;
      INIT_19             : bit_vector;
      INIT_1A             : bit_vector;
      INIT_1B             : bit_vector;
      INIT_1C             : bit_vector;
      INIT_1D             : bit_vector;
      INIT_1E             : bit_vector;
      INIT_1F             : bit_vector;
      INIT_20             : bit_vector;
      INIT_21             : bit_vector;
      INIT_22             : bit_vector;
      INIT_23             : bit_vector;
      INIT_24             : bit_vector;
      INIT_25             : bit_vector;
      INIT_26             : bit_vector;
      INIT_27             : bit_vector;
      INIT_28             : bit_vector;
      INIT_29             : bit_vector;
      INIT_2A             : bit_vector;
      INIT_2B             : bit_vector;
      INIT_2C             : bit_vector;
      INIT_2D             : bit_vector;
      INIT_2E             : bit_vector;
      INIT_2F             : bit_vector;
      INIT_30             : bit_vector;
      INIT_31             : bit_vector;
      INIT_32             : bit_vector;
      INIT_33             : bit_vector;
      INIT_34             : bit_vector;
      INIT_35             : bit_vector;
      INIT_36             : bit_vector;
      INIT_37             : bit_vector;
      INIT_38             : bit_vector;
      INIT_39             : bit_vector;
      INIT_3A             : bit_vector;
      INIT_3B             : bit_vector;
      INIT_3C             : bit_vector;
      INIT_3D             : bit_vector;
      INIT_3E             : bit_vector;
      INIT_3F             : bit_vector;
      INIT_40             : bit_vector;
      INIT_41             : bit_vector;
      INIT_42             : bit_vector;
      INIT_43             : bit_vector;
      INIT_44             : bit_vector;
      INIT_45             : bit_vector;
      INIT_46             : bit_vector;
      INIT_47             : bit_vector;
      INIT_48             : bit_vector;
      INIT_49             : bit_vector;
      INIT_4A             : bit_vector;
      INIT_4B             : bit_vector;
      INIT_4C             : bit_vector;
      INIT_4D             : bit_vector;
      INIT_4E             : bit_vector;
      INIT_4F             : bit_vector;
      INIT_50             : bit_vector;
      INIT_51             : bit_vector;
      INIT_52             : bit_vector;
      INIT_53             : bit_vector;
      INIT_54             : bit_vector;
      INIT_55             : bit_vector;
      INIT_56             : bit_vector;
      INIT_57             : bit_vector;
      INIT_58             : bit_vector;
      INIT_59             : bit_vector;
      INIT_5A             : bit_vector;
      INIT_5B             : bit_vector;
      INIT_5C             : bit_vector;
      INIT_5D             : bit_vector;
      INIT_5E             : bit_vector;
      INIT_5F             : bit_vector;
      INIT_60             : bit_vector;
      INIT_61             : bit_vector;
      INIT_62             : bit_vector;
      INIT_63             : bit_vector;
      INIT_64             : bit_vector;
      INIT_65             : bit_vector;
      INIT_66             : bit_vector;
      INIT_67             : bit_vector;
      INIT_68             : bit_vector;
      INIT_69             : bit_vector;
      INIT_6A             : bit_vector;
      INIT_6B             : bit_vector;
      INIT_6C             : bit_vector;
      INIT_6D             : bit_vector;
      INIT_6E             : bit_vector;
      INIT_6F             : bit_vector;
      INIT_70             : bit_vector;
      INIT_71             : bit_vector;
      INIT_72             : bit_vector;
      INIT_73             : bit_vector;
      INIT_74             : bit_vector;
      INIT_75             : bit_vector;
      INIT_76             : bit_vector;
      INIT_77             : bit_vector;
      INIT_78             : bit_vector;
      INIT_79             : bit_vector;
      INIT_7A             : bit_vector;
      INIT_7B             : bit_vector;
      INIT_7C             : bit_vector;
      INIT_7D             : bit_vector;
      INIT_7E             : bit_vector;
      INIT_7F             : bit_vector;
      INITP_00            : bit_vector;
      INITP_01            : bit_vector;
      INITP_02            : bit_vector;
      INITP_03            : bit_vector;
      INITP_04            : bit_vector;
      INITP_05            : bit_vector;
      INITP_06            : bit_vector;
      INITP_07            : bit_vector;
      INITP_08            : bit_vector;
      INITP_09            : bit_vector;
      INITP_0A            : bit_vector;
      INITP_0B            : bit_vector;
      INITP_0C            : bit_vector;
      INITP_0D            : bit_vector;
      INITP_0E            : bit_vector;
      INITP_0F            : bit_vector
      );
    port (
      DOA    : out std_logic_vector;
      DOB    : out std_logic_vector;
      ADDRA  : in  std_logic_vector;
      ADDRB  : in  std_logic_vector;
      CLKA   : in  std_ulogic;
      CLKB   : in  std_ulogic;
      DIA    : in  std_logic_vector;
      DIB    : in  std_logic_vector;
      ENA    : in  std_ulogic;
      ENB    : in  std_ulogic;
      REGCEA : in  std_ulogic;
      REGCEB : in  std_ulogic;
      RSTA   : in  std_ulogic;
      RSTB   : in  std_ulogic;
      WEA    : in  std_logic_vector;
      WEB    : in  std_logic_vector
      );
  end component;
end package vcomponents;
