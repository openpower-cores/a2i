-- © IBM Corp. 2020
-- Licensed under the Apache License, Version 2.0 (the "License"), as modified by
-- the terms below; you may not use the files in this repository except in
-- compliance with the License as modified.
-- You may obtain a copy of the License at http://www.apache.org/licenses/LICENSE-2.0
--
-- Modified Terms:
--
--    1) For the purpose of the patent license granted to you in Section 3 of the
--    License, the "Work" hereby includes implementations of the work of authorship
--    in physical form.
--
--    2) Notwithstanding any terms to the contrary in the License, any licenses
--    necessary for implementation of the Work that are available from OpenPOWER
--    via the Power ISA End User License Agreement (EULA) are explicitly excluded
--    hereunder, and may be obtained from OpenPOWER under the terms and conditions
--    of the EULA.  
--
-- Unless required by applicable law or agreed to in writing, the reference design
-- distributed under the License is distributed on an "AS IS" BASIS, WITHOUT
-- WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. See the License
-- for the specific language governing permissions and limitations under the License.
-- 
-- Additional rights, including the ability to physically implement a softcore that
-- is compliant with the required sections of the Power ISA Specification, are
-- available at no cost under the terms of the OpenPOWER Power ISA EULA, which can be
-- obtained (along with the Power ISA) here: https://openpowerfoundation.org. 

			

--********************************************************************
--*
--* TITLE: IU Microcode Code
--*
--* NAME: iuq_uc_rom.vhdl
--*
--*********************************************************************

library ieee,ibm,support,tri;
use ieee.std_logic_1164.all;
use ibm.std_ulogic_unsigned.all;
use ibm.std_ulogic_support.all;
use ibm.std_ulogic_function_support.all;
use support.power_logic_pkg.all;
use tri.tri_latches_pkg.all;

entity iuq_uc_rom is
  generic(ucode_width           : integer := 71;
          regmode               : integer := 6;
          expand_type           : integer := 2);
port(
     vdd                        : inout power_logic;
     gnd                        : inout power_logic;
     nclk                       : in clk_logic;
     pc_iu_func_sl_thold_0_b    : in std_ulogic;
     pc_iu_sg_0                 : in std_ulogic;
     forcee : in std_ulogic;
     d_mode                     : in std_ulogic;
     delay_lclkr                : in std_ulogic;
     mpw1_b                     : in std_ulogic;
     mpw2_b                     : in std_ulogic;
     scan_in                    : in std_ulogic;
     scan_out                   : out std_ulogic;

     rom_act                    : in std_ulogic;
     rom_addr                   : in std_ulogic_vector(0 to 9);
     rom_data                   : out std_ulogic_vector(0 to ucode_width-1)
);
-- synopsys translate_off
-- synopsys translate_on
end iuq_uc_rom;
ARCHITECTURE IUQ_UC_ROM
          OF IUQ_UC_ROM
          IS
--@@  Signal Declarations
SIGNAL ROM32_INSTR_PT                    : STD_ULOGIC_VECTOR(1 TO 893)  := 
(OTHERS=> 'U');
SIGNAL ROM64_INSTR_PT                    : STD_ULOGIC_VECTOR(1 TO 890)  := 
(OTHERS=> 'U');
SIGNAL count_src                         : STD_ULOGIC_VECTOR(0 TO 2)  := 
"UUU";
SIGNAL cr_bf2fxm                         : STD_ULOGIC  := 
'U';
SIGNAL ep                                : STD_ULOGIC  := 
'U';
SIGNAL extRT                             : STD_ULOGIC  := 
'U';
SIGNAL extS1                             : STD_ULOGIC  := 
'U';
SIGNAL extS2                             : STD_ULOGIC  := 
'U';
SIGNAL extS3                             : STD_ULOGIC  := 
'U';
SIGNAL loop_addr                         : STD_ULOGIC_VECTOR(0 TO 9)  := 
"UUUUUUUUUU";
SIGNAL loop_begin                        : STD_ULOGIC  := 
'U';
SIGNAL loop_end                          : STD_ULOGIC  := 
'U';
SIGNAL loop_init                         : STD_ULOGIC_VECTOR(0 TO 2)  := 
"UUU";
SIGNAL sel0_5                            : STD_ULOGIC  := 
'U';
SIGNAL sel11_15                          : STD_ULOGIC_VECTOR(0 TO 1)  := 
"UU";
SIGNAL sel16_20                          : STD_ULOGIC_VECTOR(0 TO 1)  := 
"UU";
SIGNAL sel21_25                          : STD_ULOGIC_VECTOR(0 TO 1)  := 
"UU";
SIGNAL sel26_30                          : STD_ULOGIC  := 
'U';
SIGNAL sel31                             : STD_ULOGIC  := 
'U';
SIGNAL sel6_10                           : STD_ULOGIC_VECTOR(0 TO 1)  := 
"UU";
SIGNAL skip_cond                         : STD_ULOGIC  := 
'U';
SIGNAL skip_zero                         : STD_ULOGIC  := 
'U';
SIGNAL template                          : STD_ULOGIC_VECTOR(0 TO 31)  := 
"UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU";
SIGNAL ucode_end                         : STD_ULOGIC  := 
'U';
SIGNAL ucode_end_early                   : STD_ULOGIC  := 
'U';
constant rom_addr_offset        : natural := 0;
constant scan_right             : natural := rom_addr_offset + 10 - 1;
-- Latches
signal rom_addr_d               : std_ulogic_vector(0 to 9);
signal rom_addr_l2              : std_ulogic_vector(0 to 9);
signal siv              : std_ulogic_vector(0 to scan_right);
signal sov              : std_ulogic_vector(0 to scan_right);
signal rom_unused       : std_ulogic;
-- synopsys translate_off
-- synopsys translate_on
  BEGIN --@@ START OF EXECUTABLE CODE FOR IUQ_UC_ROM

--64-bit core
c64: if (regmode = 6) generate
begin


-- When expanded, ROM_INSTR_PT needs more bits for 32-bit generate than 64-bit.
-- This gets rid of sourceless/sinkless warnings in 64-bit mode.
ROM32_INSTR_PT  <=  (others => '0');
rom_unused  <=  or_reduce(ROM32_INSTR_PT);
--
-- Final Table Listing
--      *INPUTS*========*OUTPUTS*===============================================================================================*
--      |               |                                                                                                       |
--      | rom_addr_l2   | template                         ucode_end                                                            |
--      | |             | |                                | ucode_end_early                                                    |
--      | |             | |                                | | loop_begin                                                       |
--      | |             | |                                | | | loop_end                                                       |
--      | |             | |                                | | | | count_src                                                    | -- Can DC if not (loop_begin or loop_end)
--      | |             | |                                | | | | |                                                            |
--      | |             | |                                | | | | |    extRT                                                   |
--      | |             | |                                | | | | |    | extS1                                                 |
--      | |             | |                                | | | | |    | | extS2                                               |
--      | |             | |                                | | | | |    | | | extS3                                             |
--      | |             | |                                | | | | |    | | | |                                                 |
--      | |             | |                                | | | | |    | | | |  sel0_5                                         |
--      | |             | |                                | | | | |    | | | |  | sel6_10                                      |
--      | |             | |                                | | | | |    | | | |  | |  sel11_15                                  |
--      | |             | |                                | | | | |    | | | |  | |  |  sel16_20                               |
--      | |             | |                                | | | | |    | | | |  | |  |  |  sel21_25                            |
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  sel26_30                         |
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | sel31                          |
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | |                              |
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | |  cr_bf2fxm                   |
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | skip_cond                 |
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | skip_zero               | -- Can DC if loop_begin not set
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | | loop_addr             | -- Can DC if loop_end not set
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | | |          loop_init  | -- 1 less than # of times to loop; Can DC if not loop_begin or not count_src=111
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | | |          |   ep     |
--      | |             | |         1111111111222222222233 | | | | |    | | | |  | |  |  |  |  | |  | | | |          |   |      |
--      | 0123456789    | 01234567890123456789012345678901 | | | | 012  | | | |  | 01 01 01 01 | |  | | | 0123456789 012 |      |
--      *TYPE*==========+=======================================================================================================+
--      | PPPPPPPPPP    | SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSS S S S S SSS  S S S S  S SS SS SS SS S S  S S S SSSSSSSSSS SSS S      |
--      *POLARITY*----->| ++++++++++++++++++++++++++++++++ + + + + +++  + + + +  + ++ ++ ++ ++ + +  + + + ++++++++++ +++ +      |
--      *PHASE*-------->| TTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTT T T T T TTT  T T T T  T TT TT TT TT T T  T T T TTTTTTTTTT TTT T      |
--      *OPTIMIZE*----->|  AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA B B B B CCC  X X X X  X XX XX XX XX X X  X X X XXXXXXXXXX XYX X       |
--      *TERMS*=========+=======================================================================================================+
--    1 | -100000000    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--    2 | -1-0000000    | .1111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--    3 | 0-11000000    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--    4 | 10-1000000    | .1...1....1.............1.1.111. . . . . ...  1 1 . .  . .. .. .1 .. . .  . . . .......... ... .      |
--    5 | 000-000000    | ..111...........111111111111111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--    6 | 110-000000    | .11111....1..........1.1111111.. . . . . ...  1 . . .  . .. .. 1. .. . .  . . . .......... ... .      |
--    7 | 011-000000    | .....1...11...1...........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--    8 | -0-0100000    | .1...1................1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--    9 | 0001100000    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   10 | 01-1100000    | .1111...........1....1........1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   11 | -01-100000    | .1.1.1...1....1......11.1.11.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   12 | -000-00000    | ................................ . . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   13 | 11-0-00000    | .........1....1.....1.11.1...... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   14 | 0001010000    | .11111....1.............1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   15 | 0-11010000    | .11111...11...11...1..1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   16 | 10-1010000    | ................................ . . . . ...  . . . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   17 | 0000110000    | .1.1......1...1.11..........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   18 | 01-0110000    | .11111.............11.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   19 | ---0110000    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   20 | 0-11110000    | ..111.....1.....1111............ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   21 | 01-1110000    | .1.1.1........1.1111111..111..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   22 | 110-110000    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   23 | 0000-10000    | ................................ . . . . ...  . . 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   24 | 1101-10000    | ................................ . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   25 | 011--10000    | .1111....1....1....1.111.11..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   26 | 11-00-0000    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   27 | 00010-0000    | ................................ . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   28 | 10-01-0000    | ..111........................1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   29 | 11011-0000    | 1..11....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   30 | 011-1-0000    | ......................1.1.1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   31 | 1-1-1-0000    | .............................1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   32 | 00--1-0000    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   33 | 1001--0000    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   34 | 101---0000    | .1.1......1...1.11..........1.1. . . . . ...  . 1 . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   35 | 111---0000    | 1..111..............1.....11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   36 | --10001000    | .1111....1....1.....1111111..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   37 | 10-1001000    | ................................ . . . . ...  . . . .  . .. 11 .. .. . .  . . . ....1111.. ... .      |
--   38 | 110-001000    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   39 | -01-001000    | ..111.....1.....11111111........ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   40 | 11-0101000    | ................................ . . . . ...  . . . .  . 11 .. .1 .. . .  . . . .......... ... .      |
--   41 | 0001101000    | .11111....1.............1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   42 | 0-11101000    | .11111...11...1....11....1.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   43 | 01-1101000    | .1111............1...11...1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   44 | 000-101000    | ................................ . . . . ...  . . 1 .  . .. .1 .. .. . .  . . . .......... ... 1      |
--   45 | 111-101000    | 1..111...11........11...1.111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   46 | 0000-01000    | ................................ . . . . ...  . . . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   47 | -11--01000    | ................................ . . . . ...  1 1 1 1  . .. .. .. .. . .  . . . .......... ... .      |
--   48 | 0001011000    | ................................ . . . . ...  1 . . .  . .. .1 .1 .1 1 .  . . . .......... ... .      |
--   49 | 0-11011000    | .1.1.1..........11111......1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   50 | 0--1011000    | ..........................1...1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   51 | 00-0111000    | .1...1....1.............1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   52 | 110-111000    | .1.1.1....1...1...........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   53 | 0-1-111000    | .11111...11...11...1..1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   54 | 0100-11000    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   55 | 1101-11000    | .1.......1....1.11............1. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   56 | 101--11000    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   57 | 011--11000    | .....1....1....1...1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   58 | -0100-1000    | .........1...........1....1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   59 | -0001-1000    | ................................ . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... 1      |
--   60 | 00-01-1000    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   61 | 10011-1000    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   62 | 11011-1000    | ................................ . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   63 | 000000-000    | ................................ . . . . ...  1 . . .  . .. .1 .. .1 1 1  . . . .......... ... .      |
--   64 | -01000-000    | .1.1.1........1.1...........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   65 | 10-000-000    | 1...1........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   66 | ---010-000    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   67 | 01-110-000    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   68 | 11-0-0-000    | .1...1....................111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   69 | 101--0-000    | .11111....................111... . . . . ...  1 . . .  . 11 .. .1 .. . .  . . . .......... ... .      |
--   70 | 000001-000    | .1.1.1...1....1..1...1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   71 | 0-1011-000    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   72 | -------000    | ................................ . . . . 1..  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   73 | 0100000100    | .11111....1...1....1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   74 | 0001000100    | 1...1.....1..................... . . . . ...  1 1 . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   75 | 1101000100    | .1.1......1...1.1...........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   76 | 0-11000100    | ...1.................11...1..11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   77 | 01-1000100    | .1111.........111111....1.....1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   78 | 011-000100    | .1111............1...11...1...1. . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   79 | 10--000100    | ..1.1..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   80 | 0100100100    | ...11.........111111....1.....1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   81 | 11-0100100    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   82 | 0001100100    | .11111....................111... . . . . ...  . . . .  . 11 .. .1 .. . .  . . . .......... ... .      |
--   83 | 0-11100100    | .1.1.1.........11....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   84 | 1-1-100100    | 1..111...11...1....1......111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   85 | 10--100100    | ................................ . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   86 | 0000-00100    | .1.1.1...1....1..1...1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   87 | 10-0-00100    | ................................ . . . . ...  . . . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   88 | 1101-00100    | ................................ . . . . ...  . . 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   89 | 0100010100    | .1111.........11111....1......1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   90 | 11-0010100    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   91 | 0001010100    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   92 | 01-1010100    | .1111.........11..........1...1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   93 | -01-010100    | .1.1.1...1....1......1111.1111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   94 | --1-010100    | ................................ . . . . ...  . 1 . 1  . .. .. .. .. . .  . . . .......... ... .      |
--   95 | 0000110100    | .11111....................111... . . . . ...  1 . . .  . 11 .. .1 .. . .  . . . .......... ... .      |
--   96 | 01-0110100    | .1111.........111....1........1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   97 | 01-1110100    | .1111....1....1...11.11..11..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   98 | 110-110100    | ..111.....1.....1111111111111..1 . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   99 | 0001-10100    | .1.1......1...1.11..........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   100 | 1101-10100    | .1...1...1.............11.1.111. . . . . ...  . 1 . 1  . .. .. .1 .. . .  . . . .......... ... .      |
--   101 | 011--10100    | .11111.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   102 | -0100-0100    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   103 | 10-01-0100    | ...............................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   104 | 11011-0100    | .1111....1....1.11............1. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   105 | 101---0100    | .1...1...1..............1.1.111. . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   106 | 0100001100    | .1111.........111111....1.....1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   107 | 0001001100    | ................................ . . . . ...  1 . . .  . 11 .. .1 .. . .  . . . .......... ... .      |
--   108 | -001001100    | .11111....................111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   109 | --11001100    | .11111.............1......11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   110 | 01-1001100    | .1111.........111.1....1......1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   111 | -1-1001100    | .................1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   112 | 00-0101100    | 1...1.....1..................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   113 | 10-0101100    | .1.1......1...1.1.....1....1111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   114 | 01-0101100    | ...11.........11111....1......1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   115 | 11-0101100    | ...1.1..................1.1.111. . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... 1      |
--   116 | 01-1101100    | .11111...11....1..........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   117 | 0-1-101100    | .1.1.1....1...1.1....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   118 | 011--01100    | .1.1.1........1.1111111..111..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   119 | 11-0011100    | 1...1....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   120 | --11011100    | ................................ . . . . ...  1 . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   121 | 01-1011100    | ...............111....1.......1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   122 | -1-1111100    | ..........1....1................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   123 | 100-111100    | ................................ . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   124 | 110-111100    | .11111...1.............11.1.111. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   125 | 0-1-111100    | ..........1...1..........1..1... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   126 | 11--111100    | ................................ . . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   127 | 0000-11100    | .1.1......1...1.11..........111. . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   128 | 0100-11100    | .....1....1...1....1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   129 | 0001-11100    | 1...1.....1..................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   130 | 11-1-11100    | ................................ . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   131 | 0-0--11100    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   132 | 011--11100    | .....1...11...1...........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   133 | 10-00-1100    | ...1.1................1....1.1.. . . . . ...  1 . . .  . .. .1 .1 .. . .  . . . .......... ... .      |
--   134 | -1110-1100    | 1........................1..11.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   135 | 1-1-0-1100    | ................................ . . . . ...  1 . . 1  . .. 1. 11 .. . .  . . . .......... ... .      |
--   136 | 00011-1100    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   137 | 1-011-1100    | .1...1...1.............11.1.111. . . . . ...  . 1 . .  . .. .. .1 .. . .  . . . .......... ... 1      |
--   138 | -01-00-100    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   139 | 11-010-100    | ....1.....1...1................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   140 | 101--0-100    | .11111....1.............1.1.111. . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   141 | 000001-100    | ................................ . . . . ...  1 . . .  . .. .1 .1 .1 1 1  . . . .......... ... .      |
--   142 | 00-001-100    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   143 | 1-1-01-100    | 1...11...11.............11111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   144 | -00111-100    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   145 | 0-1111-100    | .11111.............1......11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   146 | 10-0-1-100    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   147 | 11-0000-00    | ..111..........................1 . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   148 | -010100-00    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   149 | ---0100-00    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   150 | -010010-00    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   151 | 10--010-00    | ..111........................... . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   152 | --1---0-00    | ................................ . . . . ...  1 . 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   153 | 0000001-00    | .11111....1.............1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   154 | -010001-00    | .........1...........1....1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   155 | 10-1001-00    | ...111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   156 | ----001-00    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   157 | 01-1111-00    | .....1.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   158 | 11-1111-00    | 1...11.........1........111111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   159 | -11-111-00    | ................................ . . . . ...  1 1 . 1  . .. .. .1 .. . .  . . . .......... ... .      |
--   160 | 1001-11-00    | 1..11....1.....................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   161 | 01---11-00    | .1111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   162 | 011-1-1-00    | .1...1.........1....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   163 | --0-10--00    | ................................ . . . . ...  1 . . 1  . .. .. .. .. . .  . . . ......1... ... .      |
--   164 | 10-001--00    | .1.1.1................1....1.1.. . . . . ...  1 . . .  . .. .1 .1 .. . .  . . . .......... ... .      |
--   165 | --10-1--00    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   166 | 1101-1--00    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   167 | 0-1-1---00    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   168 | 0100000010    | ..1111....1....1.1.1.1.1.1.1.1.1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   169 | 1101000010    | .1.1.1....1...1...........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   170 | 0-11000010    | .1...1.........1........11.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   171 | 10-1000010    | .1.1......1...1.1.....1....1111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   172 | 011-000010    | .1111....1....1...1..11.111..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   173 | 11-0100010    | .1111.....1....1.1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   174 | 0-11100010    | ..111....11...11..........1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   175 | 01-1100010    | .1111..........111....1.......1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   176 | 0000-00010    | 1...1....1.....................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   177 | 1-1--00010    | 1..111...1................11..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   178 | -0---00010    | ................................ . . . . ...  . . 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   179 | -010010010    | 1..11....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   180 | 00-1110010    | .1.1.1...1....1......111.1111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   181 | 01-1110010    | ...111...11...1...........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   182 | 110-110010    | ...11..............1.1...1.1.... . . . . ...  . . 1 .  . .1 .. .. .. . .  . . . .......... ... .      |
--   183 | -11-110010    | 1..111...11...............11..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   184 | 0100-10010    | .1111.....1...1......11111...11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   185 | 11-0-10010    | .1...1....1.............1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   186 | 0001-10010    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   187 | 1101-10010    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   188 | 011--10010    | .1111...........11...11...1...1. . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   189 | 11-00-0010    | ................................ . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   190 | 1--00-0010    | ..1............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   191 | 0-110-0010    | ..111.....1.....11.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   192 | 1-1-0-0010    | ................................ . . . . ...  1 . . 1  . .. .1 .. .. . .  . . . .......... ... .      |
--   193 | 00011-0010    | .11.1....1...................... . . . . ...  . 1 . .  . .. 11 .. .. . .  . . . .......... ... .      |
--   194 | 11011-0010    | ...111....1..........1.11111111. . . . . ...  . . . .  . .. .. 1. .. . .  . . . .......... ... .      |
--   195 | 1--11-0010    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   196 | 011-1-0010    | .1...1........1.....1.1..1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   197 | 111-1-0010    | ................................ . . . . ...  . . . .  . .. .. .. 1. . .  . . . .......... ... .      |
--   198 | 101---0010    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   199 | 1--0001010    | .1.1......1...1.11..........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   200 | 1101001010    | ................................ 1 . . . ...  . . . .  . 1. .1 .1 .1 1 1  . . . .......... ... .      |
--   201 | 00-1001010    | .1.1.1...1....1......111..111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   202 | 0-0-001010    | .1111.....1...1......11111...11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   203 | 011-001010    | .11111....1....1...1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   204 | 10--001010    | .....1....1.............1.1.111. . . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   205 | 0-11101010    | .11111.............1.1....11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   206 | 01-1101010    | .11111.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   207 | 110-101010    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   208 | 0001-01010    | .1111....1....1.11............1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   209 | 1-01-01010    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   210 | 000--01010    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   211 | 11-0011010    | ...111.........1......1....1.1.. . . . . ...  . 1 1 .  . 1. .. .. .. . .  . . . .......... ... .      |
--   212 | 1--0011010    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   213 | --11011010    | .........11...11..............1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   214 | 01-1011010    | .1.............11....1........1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   215 | -0-0111010    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   216 | 01-1111010    | .1111....1....1.....1111111..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   217 | 1-0-111010    | .1.1......1...1.1...........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   218 | 0-1-111010    | .1.1.1.........11..1..111.11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   219 | 0100-11010    | ..1111....1....1.1.1.1.1.1.1.1.1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   220 | -010-11010    | ................................ . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   221 | 1001-11010    | 1..11....1....................1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   222 | 1101-11010    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   223 | 011--11010    | .1.1.1........1.1111111..111..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   224 | 00010-1010    | ...............................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   225 | -0101-1010    | 1..11....1...................... . . . . ...  . 1 . 1  . .. .. .1 .1 1 .  . . . .......... ... .      |
--   226 | 10-01-1010    | .1.1.1...1....1.11........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   227 | -0-1--1010    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   228 | 000100-010    | ..111..........................1 . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   229 | 01-100-010    | .1111.....1...1......11111...11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   230 | 010010-010    | .1111.....1...1......11111...11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   231 | 101--0-010    | ..111..........................1 . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   232 | 000001-010    | ................................ . . . . ...  . 1 . .  . .. 11 .. .. . .  . . . .......... ... .      |
--   233 | 1-1-01-010    | 1..111....................11..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   234 | --1011-010    | ................................ . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   235 | --01-1-010    | ................................ . . . . ...  1 1 . 1  . .. .. .. .. . .  . . . 1....1.... 1.. .      |
--   236 | 0100000110    | ...............1...11........... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   237 | 11-0000110    | 1...1.....1..................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   238 | 0001000110    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   239 | 1101000110    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   240 | --11000110    | ..111....11...11...........1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   241 | 10-1000110    | .1...1....1.............1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   242 | 11-1000110    | 1..11....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   243 | 010-000110    | .11111...1................111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   244 | 011-000110    | .1...1.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   245 | 0000100110    | ...1.1...1...........111..11.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   246 | 0001100110    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   247 | 0-01100110    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   248 | 0000-00110    | ................................ . . . . ...  . . . .  . .. 1. .. .. . .  . . . .......... ... .      |
--   249 | 0100-00110    | ...1.1...1................111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   250 | -010-00110    | ................................ . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   251 | 10-1-00110    | ................................ . . . . ...  . . . 1  . .. .. .1 .. . .  . . . .......... ... .      |
--   252 | 11-0010110    | .1.1......1...1.11..........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   253 | 0001010110    | ..111.....1.....11111111111111.1 . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   254 | 0-11010110    | .11111.............1......11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   255 | -000110110    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   256 | --01110110    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   257 | 01-1110110    | .1111...........11...11...1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   258 | 110-110110    | .11111....1..........1.11.111.1. . . . . ...  1 . . .  . .. .. 1. .. . .  . . . .......... ... .      |
--   259 | 1001-10110    | 1..11....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   260 | 1101-10110    | .11111....1..........1.11111111. . . . . ...  . . . .  . .. .. 1. .. . .  . . . .......... ... .      |
--   261 | 011--10110    | .1111....1....1.....1111111..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   262 | 1-1-0-0110    | .........1.........11...1....... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   263 | 10011-0110    | .1...1...1.............11.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   264 | 0-111-0110    | .1.1.1....1...1.1....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   265 | -100001110    | .11111...1................111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   266 | -010001110    | ................................ . . . . ...  1 . . .  . .. .1 .1 .1 1 1  . . . .......... ... .      |
--   267 | 11-0001110    | ................................ . . . . ...  1 . . .  . 11 .. .1 .. . .  . . . .......... ... .      |
--   268 | 0-11001110    | .1.1.1....1...1.1....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   269 | 01-1001110    | .11111.............1......111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   270 | 0000101110    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   271 | 10-0101110    | .1.1......1...1..1...1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   272 | 0-11101110    | ...1.1....1...11...1..1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   273 | -1-1101110    | .1111.....1....1..11111...1..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   274 | 11--101110    | ...11....1....1.11............1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   275 | 1101-01110    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   276 | 011--01110    | .1...1...11...1...........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   277 | 11-0011110    | .1111....1....1..1...1.1111..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   278 | --11011110    | .....1....1....1........11.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   279 | -01-011110    | ................................ . . . . ...  1 1 . 1  . .. .. .1 .. . .  . . . .......... ... 1      |
--   280 | -1-1111110    | .1.1.1........1.1111111..111..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   281 | -0--111110    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   282 | 11--111110    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   283 | 0000-11110    | ..........1.....11111111111111.. . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   284 | 0100-11110    | .11111...1.....1...11.....111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   285 | -010-11110    | .1...1...1.............11.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   286 | 0001-11110    | .1.......1....1.11............1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   287 | 10-1-11110    | .1.1.1........1..1........1111.. . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   288 | 11-1-11110    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   289 | -1---11110    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . 11..1111.. ... .      |
--   290 | 01-01-1110    | ...111.............1......111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   291 | 00011-1110    | ................................ . . . . ...  . 1 . .  . .. 11 .. .. . .  . . . .......... ... .      |
--   292 | 00-11-1110    | .11.1....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   293 | 1--11-1110    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   294 | 111-10-110    | 1..111........11........111111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   295 | --10-0-110    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   296 | 000001-110    | 1..............................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   297 | 0-1011-110    | .1...1...1.............11.1.111. . . . . ...  . 1 . 1  . .. .. .1 .. . .  . . . .......... ... 1      |
--   298 | -00111-110    | .1.1..........1......11...11111. . . . . ...  . . 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   299 | 11011--110    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   300 | -1111--110    | ................................ . . . . ...  1 1 . 1  . .. .. .1 .. . .  . . . .......... ... .      |
--   301 | 10--1--110    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . 1 1...1..1.1 ... .      |
--   302 | 101----110    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   303 | -010000-10    | ................................ . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   304 | 0000110-10    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   305 | 10-0110-10    | .1.1.1...1....1..1........1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   306 | 100-110-10    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   307 | --101-0-10    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   308 | 0000001-10    | .1...1.............11...1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   309 | 000-001-10    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   310 | 11-0101-10    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   311 | 111-101-10    | 1..111...1....11........111111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   312 | 0000011-10    | .....1...............111..11.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   313 | 00--011-10    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   314 | -001111-10    | ...............................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   315 | 101--11-10    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   316 | 00010-1-10    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   317 | -0-100--10    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . 1..1..11.1 ... .      |
--   318 | 01---0--10    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   319 | 1-0111--10    | ...111...1.............11.1.111. . . . . ...  . . . .  . .. .. .1 .. . .  . . 1 .......... ... .      |
--   320 | 00000---10    | ....1....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   321 | 1--00000-0    | ................................ . . . . ...  . . . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   322 | -0101000-0    | .1.......1....1.11............1. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   323 | 10-0-000-0    | ................................ . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   324 | 10-10100-0    | ..111........................1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   325 | 01-10100-0    | .11111.............11.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   326 | -01-0100-0    | ................................ . . . . ...  . 1 . 1  . .. .. .. .. . .  . . . .......... ... .      |
--   327 | 11-00-00-0    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   328 | 1-011-00-0    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . 1..11..1.1 ... .      |
--   329 | -0-00010-0    | .................1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   330 | 11-00010-0    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   331 | 000-0010-0    | .1.1......1...1.11..........111. . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   332 | 0000-010-0    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   333 | 1--00110-0    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   334 | 0-010110-0    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   335 | 110-1110-0    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   336 | 10-000-0-0    | ................................ . . . . ...  . . . .  . .1 .. .1 .. . .  . . . .......... ... .      |
--   337 | --110001-0    | ................................ . . . . ...  1 1 1 1  . .. .. .. .. . .  . . . .......... ... .      |
--   338 | -10-0001-0    | ................................ . . . . ...  1 1 . 1  . .. .. .. .. . .  . . . .......... ... .      |
--   339 | 1-1-0001-0    | 1..111....1..............1111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   340 | 10-01001-0    | ..111........................1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   341 | 01-11001-0    | ..111....1.....................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   342 | 10-1-001-0    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   343 | -0100101-0    | .................1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   344 | 11-00101-0    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   345 | 11-0-011-0    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   346 | 1--11111-0    | ................................ . . . . ...  . . 1 .  . .1 .. .. .. . .  . . . .......... ... .      |
--   347 | 10-1-111-0    | ..............................1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   348 | 101--111-0    | ...111.............1.1..11111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   349 | 0-101-11-0    | .1.......1....1.11............1. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   350 | -1111-11-0    | 1..111.........1..........1...1. . . . . ...  . 1 1 1  . .1 .. .. .. . 1  . . . .......... ... .      |
--   351 | -1-010-1-0    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   352 | -01011-1-0    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   353 | 011-1--1-0    | ...111.........1....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   354 | 10-0000--0    | 1............................... . . . . ...  . . . .  . .1 .1 .1 .1 1 1  . . . .......... ... .      |
--   355 | -110110--0    | 1....1...1................1..... . . . . ...  1 . . .  . .. .. 11 .. . .  . . . .......... ... .      |
--   356 | 0000001--0    | ................................ . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... 1      |
--   357 | 10--001--0    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   358 | 1-1-011--0    | 1...11.........1..........1...1. . . . . ...  . 1 1 1  . .1 .. .. .. . 1  . . . .......... ... .      |
--   359 | -001111--0    | 1..11....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   360 | 10-00-1--0    | ....1........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   361 | -100000001    | ..111.....1......1.1.1.1.1.1.1.1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   362 | 0001000001    | 1...1....1...................... . . . . ...  . . . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   363 | 0-11000001    | ...............11....1.......... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   364 | 110-000001    | .1.1.1....1...1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   365 | 011-000001    | .1111....1....1.....1111111..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   366 | 0-11100001    | .11111...11...1.........11.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   367 | 1-1-100001    | 1....1....1...............11..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   368 | 0000-00001    | 1...1.....1..................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   369 | 11-0-00001    | .1111....1....1.11............1. . . 1 . ...  . . . .  . .. .. .. .. . .  . 1 . .......... 1.. .      |
--   370 | 01-0010001    | .....1.........1................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   371 | 01-1010001    | .1111.........111....1........1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   372 | 000-010001    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   373 | -000110001    | ................................ . . . . ...  . 1 1 .  . .. 11 .. .. . .  . . . 1...1.1..1 ... .      |
--   374 | 01-0110001    | ..111.....1...............111111 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   375 | 00-1110001    | .1.1.1....1...1.1....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   376 | -00-110001    | ................................ . 1 . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   377 | 110-110001    | .11.1.....1...1................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   378 | -11-110001    | 1..111....................11..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   379 | 1101-10001    | .11111...1.............11.1.111. . . 1 . ...  . 1 . 1  . .. .. .1 .. . .  . . . .......... ... .      |
--   380 | 10-1-10001    | ................................ . . . . ...  . . 1 .  . .1 .. .. .. . .  . . . .......... ... .      |
--   381 | 011--10001    | .1111.....1........1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   382 | 1-1--10001    | .........1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   383 | 11-00-0001    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   384 | 1-1-0-0001    | 1..111....1...............1111.. . . . . ...  1 . 1 1  . .. 1. .. .. . .  . . . .......... ... .      |
--   385 | 10011-0001    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   386 | 11011-0001    | ................................ 1 . . . ...  . . . .  . 1. .1 .. .. . .  . . . .......... ... .      |
--   387 | 101---0001    | ...................1.1..11...... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   388 | --10001001    | .1111....1....1....11111..1..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   389 | 11-1001001    | 1..11....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   390 | ---1001001    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   391 | -01-001001    | .1.1.1....1...1.1....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   392 | -000101001    | 1...1....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   393 | -0-0101001    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . 1 ..1......1 ... .      |
--   394 | 11-0101001    | .11111...1..............1.1.111. . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... 1      |
--   395 | 0001101001    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   396 | 0-11101001    | ..111....11...11...........1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   397 | 01-1101001    | .1.1.1........1.1111111..111..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   398 | 11-1101001    | ................................ . . . . ...  1 1 . 1  . .. .. .1 .. . .  . . . .......... 1.. 1      |
--   399 | 0100-01001    | .....1.........1................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   400 | 0----01001    | ................................ . . . . ...  . 1 1 .  . .. .. .. .. . .  . . . ....1..11. ... .      |
--   401 | 11-0011001    | ..111.....1.....11111111111111.1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   402 | 0001011001    | 1...1....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   403 | 01-1111001    | .11111...11...1...........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   404 | 1-0-111001    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   405 | 0000-11001    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   406 | 0100-11001    | ..111.....1......1.1.1.1.1.1.1.1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   407 | --10-11001    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   408 | 1101-11001    | .1111.....1....1.1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   409 | 0-11-11001    | .11111.............1......11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   410 | 101--11001    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   411 | 10-01-1001    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   412 | 11011-1001    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   413 | 1-011-1001    | .11111...1.............11.1.111. . . . . ...  . . . 1  . .. .. .1 .. . .  . . . .......... ... .      |
--   414 | -01000-001    | .1.1..........1......11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   415 | 11-000-001    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   416 | 01-100-001    | .....1.........1................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   417 | 01-010-001    | .....1.........1................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   418 | 101--0-001    | .11111...1..............1.1.111. . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   419 | 0-1101-001    | .11111.............1......11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   420 | 0-1011-001    | .1111.....1...1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   421 | 00--11-001    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . ....11.11. ... .      |
--   422 | 0100000101    | .1111.........1111111....1....1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   423 | 1101000101    | ................................ . . . . ...  1 . . .  . .. .1 .1 .1 1 1  . . . .......... ... .      |
--   424 | 10-1000101    | .1.1......1...1..1...1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   425 | 01-1000101    | .11111...1.....1...11.....111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   426 | 000-000101    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   427 | 011-000101    | .1.1.1........1.1111111..111..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   428 | 1-1-000101    | 1..111..................1.1111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   429 | 0100100101    | .11111...1.....1...11.....111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   430 | 11-0100101    | .11111.............1.1..1111111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   431 | 1--0100101    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   432 | 0001100101    | .1...1..................1.1.111. . . . . ...  . . 1 .  . .. .1 .. .. . .  . . . .......... ... 1      |
--   433 | 0-11100101    | .1...1.........1........11.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   434 | 01-1100101    | .1.......1....1......11111...11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   435 | 1-1-100101    | 1....1...1.....1....1.....111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   436 | 10--100101    | ................................ . . 1 . ...  . . . .  . .1 .. .. .. . .  . . 1 .......... ... .      |
--   437 | 11-0010101    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   438 | 0001010101    | .11111...1...........1111.11.1.. . . . . ...  . 1 . .  . .. 11 .. .. . .  . . . .......... ... .      |
--   439 | -101010101    | .11111.............11.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   440 | -01-010101    | .11111...11...11...1..1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   441 | 0000110101    | ...1.1..................1.1.111. . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... 1      |
--   442 | 01-1110101    | ..........1....1................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   443 | 110-110101    | .11111.........1......1....1.1.. 1 . . . ...  . . . .  . 1. .. .. .. . .  . . . .......... ... .      |
--   444 | 1101-10101    | ................................ 1 . . . ...  . . . .  . 1. .1 .1 .. . .  . . . .......... ... .      |
--   445 | 011--10101    | .11111...11...1...........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   446 | -0100-0101    | .11111...1.............11.1.111. . . . . ...  . 1 . 1  . .. .. .1 .. . .  . . . .......... ... 1      |
--   447 | 1-1-0-0101    | ................................ . . . . ...  1 . . 1  . .. 1. 11 .. . .  . . . .......... ... .      |
--   448 | 0-111-0101    | ..111.....1.....11.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   449 | --1-1-0101    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . ..1.11..11 ... .      |
--   450 | 101---0101    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   451 | 0100001101    | .11111...1.....1...11.....111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   452 | 11-0001101    | ................................ 1 . . . ...  . . . .  . 1. .1 .1 .1 1 1  . . . .......... ... .      |
--   453 | 0001001101    | .11111...1..............1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   454 | 01-1001101    | .11111.............11.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   455 | 01-0101101    | .11111.............11.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   456 | 11-0101101    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   457 | 0-11101101    | .1.1.1...1....1......111..111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   458 | 01-1101101    | .1111.....1....1....1111111..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   459 | -010-01101    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   460 | 011--01101    | .11111.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   461 | --11011101    | ...............1..........1...1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   462 | 11--011101    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   463 | -1-1111101    | .1111................11...1...1. . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   464 | 1-0-111101    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   465 | 0000-11101    | ................................ . . . . ...  . 1 . .  . .. 11 .. .. . .  . . . .......... ... .      |
--   466 | 0100-11101    | .1111.........1111111....1....1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   467 | 0001-11101    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   468 | 1001-11101    | ..111........................1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   469 | -0-1-11101    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   470 | 11-1-11101    | 1..11....1...................... . . . . ...  . . . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   471 | 11-00-1101    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   472 | 0-1100-101    | ..111.....1.....1111............ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   473 | 000010-101    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   474 | 000110-101    | ..111....1.....1................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   475 | 101--0-101    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   476 | 01---0-101    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   477 | -00001-101    | 1...1.....1..................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   478 | -01001-101    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   479 | -1001--101    | ................................ . . . . ...  . 1 1 .  . .. .. .. .. . .  . . . 11..1...1. ... .      |
--   480 | 11011--101    | .1........1....1.1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   481 | 011-1--101    | .1.1.1....1.....11....1...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   482 | 11-0000-01    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   483 | -010100-01    | .1111.....1...1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   484 | 10-1100-01    | .1.1.1........1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   485 | -010010-01    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   486 | 0--0010-01    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . ..1...1111 ... .      |
--   487 | 10-1010-01    | ................................ . . 1 . ...  1 . . .  . .1 .. .. .. . .  . . 1 .......... ... .      |
--   488 | 10-0110-01    | ...1.1........1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   489 | 0001110-01    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   490 | 01-1110-01    | .11111.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   491 | 0000001-01    | ..111....11....................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   492 | 0001001-01    | ................................ . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   493 | 10-1001-01    | .1.1.1...1....1..1........1.111. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   494 | -1-0-01-01    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   495 | -001111-01    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   496 | 100-111-01    | .....1..................1.1.111. . . 1 . ...  1 . . .  . .. .. .1 .. . .  . . 1 .......... ... .      |
--   497 | 011--11-01    | .1111................11...1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   498 | -0101-1-01    | .1111....1....1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   499 | -00011--01    | .11.1....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   500 | 00000---01    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   501 | -0011---01    | ................................ . . . . ...  1 . . .  . .. .. .. .. . .  . . . ...1...... ... .      |
--   502 | 0-------01    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   503 | 0100000011    | .1111.....1...1......11111...11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   504 | -010000011    | .1...1...1.............11.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   505 | 1101000011    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   506 | 011-000011    | .11111....1....1...1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   507 | 1-1-000011    | .........11.........1....1..1... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   508 | -010100011    | .1111.....1....1.1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   509 | 1--0100011    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   510 | 0-11100011    | .11111.............1.1....11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   511 | 0000-00011    | .1.1......1...1..1...1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   512 | 10-1-00011    | .1...1....1.............1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   513 | 10---00011    | ................................ . . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   514 | --00010011    | .11..1................1....1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   515 | -010010011    | ................................ . . . . ...  . . . .  . .. .. .. .1 1 .  . . . .......... ... .      |
--   516 | -0-0010011    | ..111........................1.. 1 . . . ...  . . 1 .  . 1. .1 .. .. . .  . . . .......... ... .      |
--   517 | 1--0010011    | ...11....1....1.....1..1.11.1... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   518 | 10--010011    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   519 | 00-1110011    | .11111...11...11...1..1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   520 | 01-1110011    | ...11....1....1.....1111111..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   521 | 0001-10011    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   522 | 1101-10011    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   523 | 011--10011    | .1.1.1........1.1111111..111..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   524 | -0100-0011    | ................................ . . . . ...  . . . 1  . .. .1 .1 .. . .  . . . .......... ... 1      |
--   525 | 0-110-0011    | .1.1.1....1...1.1....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   526 | 11--0-0011    | ................................ . . . . ...  1 1 1 1  . .. .. .. .. . .  . . . 11...1.... ... .      |
--   527 | 10-01-0011    | 1...1.....1..................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   528 | 00011-0011    | ................................ 1 . . . ...  . . . .  . 1. .1 .1 .1 1 .  . . . .......... ... .      |
--   529 | 101---0011    | ................................ . . . . ...  . . . .  . 11 .. .1 .. . .  . . . .......... ... .      |
--   530 | 1--0001011    | .1...1.............1.1..111111.. . . . . ...  . . 1 .  . .1 .. .. .. . .  . . . .......... ... .      |
--   531 | 1101001011    | .1...1....1..........1.1111111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   532 | 00-1001011    | .11111...11...11...1..1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   533 | 11-1001011    | ................................ . . . . ...  . . . .  . .. .. 1. .. . .  . . . .......... ... .      |
--   534 | 0000101011    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   535 | 11-0101011    | .1.......1....1..1...1.1111..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   536 | -001101011    | .1...............1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   537 | 01-1101011    | .1............11................ . . . . ...  . . . .  . 1. .. .. .. . .  . . . .......... ... .      |
--   538 | 0-1-101011    | ..111.....1.....11111111........ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   539 | 0100-01011    | .1...1....1...1....1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   540 | 011--01011    | .1..............1....11...1...1. . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   541 | 1--0011011    | ................................ . . . . ...  . . . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   542 | --11011011    | .11111........1....11....1.1.... 1 . . . ...  . . 1 .  . 1. .. .. .. . 1  . . . .......... ... .      |
--   543 | 0---011011    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   544 | -1-1111011    | .1.......1....1...1.111.1.1..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   545 | 0100-11011    | .1........1...1......11111...11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   546 | -010-11011    | .11111...1.............11.1.111. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   547 | 11-0-11011    | ................................ . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   548 | 11-1-11011    | .1........1...1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   549 | 00010-1011    | .1111....1....1..1...1.1111..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   550 | --101-1011    | ................................ 1 . . . ...  . . . .  . 1. .1 .1 .1 1 .  . . . .......... ... .      |
--   551 | -1----1011    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   552 | 000100-011    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   553 | 01-100-011    | .11111....1...1....1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   554 | 010010-011    | .11111....1...1....1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   555 | 10-110-011    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   556 | -00001-011    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   557 | 1-1-01-011    | 1...11....1.............11111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   558 | 000011-011    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   559 | --1011-011    | .11111...1.............11.1.111. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   560 | 000111-011    | ................................ 1 . . . ...  . . . .  . 1. .1 .1 .1 1 1  . . . .......... ... .      |
--   561 | -010-1-011    | ................................ . . . . ...  . . . 1  . .. .. .1 .. . 1  . . . .......... ... 1      |
--   562 | 00011--011    | ..111.....1....1................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   563 | 011-1--011    | .1.1.1....1.....111....1..11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   564 | 111-1--011    | 1..111.........1....1...1.1111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   565 | -1-1---011    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   566 | -010000111    | .11111................1....1.1.. . . . . ...  . 1 . .  . 1. .. .1 .. . .  . . . .......... ... .      |
--   567 | -0-0000111    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   568 | 11-0000111    | .1...1...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   569 | 0001000111    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   570 | 0-11000111    | .11111.............1.1....11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   571 | 011-000111    | .11111...11...1...........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   572 | -010100111    | 1..11....1...................... . . 1 . ...  . . . 1  . .. .. .1 .1 1 .  . . . .......... 1.. .      |
--   573 | 11-0100111    | ................................ . . . . ...  . . . .  . 1. .1 .1 .1 1 1  . . . .......... ... .      |
--   574 | 1--0100111    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   575 | 0001100111    | .1111....1....1..1...1.1111..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   576 | 0-11100111    | .1.1.1...1....1......11.1111.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   577 | 01-1100111    | .1...1.............1......111... 1 . . . ...  . 1 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   578 | -000-00111    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   579 | 0-00010111    | .1.1......1...1..1...1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   580 | 1--0010111    | .11111.............1.1..111111.. . . . . ...  . . 1 .  . .1 .. .. .. . .  . . . .......... ... .      |
--   581 | 0-01010111    | .11111.........1......1....1.1.. 1 . . . ...  . 1 1 .  . 1. .. .. .. . .  . . . .......... ... .      |
--   582 | 0-11010111    | .1.1.1.........11..1..111.11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   583 | 110-110111    | .1.1.1....1...1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   584 | 010--10111    | .1.1.1........1.1111111..111..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   585 | 01000-0111    | ...1.1.........1.........1.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   586 | 01-10-0111    | .11111..............1.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   587 | 01001-0111    | ...1.1..............1.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   588 | -000001111    | .1.1......1...1..1...1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   589 | 0100001111    | .11111..............1.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   590 | -010001111    | 1..11....1...................... . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   591 | 1--0001111    | .1...1...1..............1.1.111. . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   592 | --11001111    | .1.1.1...1....1......111.1111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   593 | 10--001111    | .11.1....1...................... 1 . . . ...  . 1 . .  . .. 11 .. .. . .  . . . .......... ... .      |
--   594 | 0---001111    | ................................ . . . . ...  1 1 . 1  . .. .. .. .. . .  . . . .......... ... .      |
--   595 | 0000101111    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   596 | 01-0101111    | .1111.........1111....1.......1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   597 | 0001101111    | ..111.....1.....1111111111111..1 . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   598 | -1-1101111    | .1111...........1....11...1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   599 | 11--101111    | .1........1....1.1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   600 | 11-1-01111    | .1.1......1...1.1...........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   601 | -0-0011111    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   602 | 1--0011111    | 1...1.....1..................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   603 | 0-01011111    | .1111.....1....1.1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   604 | 00-0111111    | .11111.........1......1....1.1.. 1 . . . ...  . 1 1 .  . 1. .. .. .. . .  . . . .......... ... .      |
--   605 | -0-1111111    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   606 | 11--111111    | .11111...1.............11.1.111. 1 . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   607 | --10-11111    | .1...1................1....1.1.. 1 . . . ...  . . . .  . 1. .1 .1 .. . .  . . . .......... ... .      |
--   608 | 10-0-11111    | .1.1.1...1....1.11........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   609 | --11-11111    | ..........1...1...........1...1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   610 | 10-1-11111    | 1..11....1...................... . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   611 | 01-1-11111    | .11111.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   612 | 11-1-11111    | .1111....1....1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   613 | 01-10-1111    | .1111.........1111....1.......1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   614 | --101-1111    | .1111.....1....1.1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   615 | 1-011-1111    | .11111...1.............11.1.111. . . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   616 | 0-111-1111    | .11111.............1......11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   617 | -11---1111    | .1111....1....1.....1111111..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   618 | 1-1---1111    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   619 | 111-10-111    | 1....1....1........11...1.111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   620 | 11-0-0-111    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   621 | 0-1011-111    | ................................ . . . . ...  . . . .  . 1. .1 .1 .. . .  . . . .......... ... .      |
--   622 | --1011-111    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   623 | 0-1111-111    | .1.1.....1....1......1.11.1.1... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   624 | -10-11-111    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   625 | 0-1-11-111    | .....1................1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   626 | 0100-1-111    | .11111.........1.........1.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   627 | 101--1-111    | .11111....1.............1.1.111. . . . . ...  . . 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   628 | 011--1-111    | .1111....1....1.....11111.1..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   629 | 011-1--111    | .1.1.1....1.....1....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   630 | -1--000-11    | ................................ . . . . ...  1 1 . 1  . .. .. .. .. . .  . . . .......... ... .      |
--   631 | --1-100-11    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   632 | 01-1010-11    | ..111.....1..............1111111 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   633 | 0000110-11    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   634 | 0001110-11    | ................................ . . . . ...  . . . .  . .. .1 .1 .1 1 1  . . . .......... ... .      |
--   635 | -001110-11    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   636 | 0100-10-11    | ...111....1...1....1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   637 | 11011-0-11    | .1........1...1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   638 | -1-0--0-11    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   639 | 0001001-11    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   640 | 01-1101-11    | ................................ . . . . ...  1 . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   641 | 10-0-01-11    | ....1.....1....................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   642 | 0-1-111-11    | .1.1.1....1...1.11111....111111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   643 | -11--11-11    | .1...1.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   644 | 1-1--11-11    | .1.1......1...1.11..........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   645 | -1110-1-11    | .........1..............1....... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   646 | 11011-1-11    | .1.......1....1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   647 | -1-1--1-11    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   648 | 11-111--11    | ................................ . . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   649 | -11-11--11    | ..............1..........1...... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   650 | -1--11--11    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   651 | 10---1--11    | ................................ . . . . ...  1 . . .  . .. .. .. .. . .  . . . .......1.. ... .      |
--   652 | 1-10----11    | ................................ . . . . ...  . 1 1 .  1 .1 .. .. .1 1 1  . . . .......... ... .      |
--   653 | 11-00000-1    | 1...1....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   654 | 10--0000-1    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   655 | 01-11000-1    | .1...1....1...........1..1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   656 | ---11000-1    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   657 | 10-10100-1    | 1..1............................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   658 | 10--0100-1    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   659 | 00011-00-1    | ..111....1.....1................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   660 | 101---00-1    | .11111....................111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   661 | -0000010-1    | ................................ . . . . ...  . . . .  . 1. .. .1 .. . .  . . . .......... ... .      |
--   662 | -0100010-1    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   663 | 00010010-1    | .11111...1...........1111.11.1.. 1 . . . ...  . . . .  . .. 1. .. .. . .  . . . .......... ... .      |
--   664 | 111-1010-1    | 1..111.........1.........11111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   665 | 11-00110-1    | ................................ . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   666 | 1001-110-1    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   667 | 101--110-1    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   668 | 10-000-0-1    | ..111........................... 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   669 | --0100-0-1    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   670 | 1--100-0-1    | ................................ . . . . ...  1 . . 1  . .. .. .. .. . .  . . . .......... ... .      |
--   671 | 0-0010-0-1    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   672 | -00101-0-1    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . ...1..111. ... .      |
--   673 | 0-1-11-0-1    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... 1.. .      |
--   674 | -1-00001-1    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . 11.....1.. ... .      |
--   675 | 11010001-1    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   676 | --1-0001-1    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   677 | -0100101-1    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   678 | 10-10101-1    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   679 | 100-1101-1    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   680 | 1-0-1101-1    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   681 | 0100-101-1    | .11111.............11.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   682 | 1101-101-1    | .1111.....1...1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   683 | 0--10-01-1    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   684 | 11010011-1    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   685 | 10-01011-1    | ....1.....1...................1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   686 | -----011-1    | ................................ . . . . ..1  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   687 | 10-00111-1    | .11...........................1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   688 | ---10111-1    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . ...1.1.... ... .      |
--   689 | ---01111-1    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   690 | 1--11111-1    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   691 | 0-1-1111-1    | ..111....11...11..............1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   692 | 1-0--111-1    | ................................ . . . . ...  . 1 . 1  . .. .. .. .. . .  . . . 1......1.1 1.. .      |
--   693 | -11--111-1    | .........1....1.....1..111...... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   694 | 10-00-11-1    | 1...1........................... . . . . ...  . 1 . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   695 | -1110-11-1    | 1..111.........1..........1...1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   696 | 0-0-0-11-1    | ................................ . . . . ...  1 . 1 .  . .. .. .. .. . .  . . . ......1.1. ... .      |
--   697 | 1-1-0-11-1    | ................................ . . . . ...  . 1 1 1  . .1 .. .. .. . 1  . . . .......... ... .      |
--   698 | 11011-11-1    | .....1................1....1.1.. . . . . ...  . . . .  . 1. .1 .1 .. . .  . . . .......... ... .      |
--   699 | 11-11-11-1    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   700 | -011-0-1-1    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . 1.111.1.1. ... .      |
--   701 | 1-1--0-1-1    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   702 | 1-1-01-1-1    | 1...11...................11111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   703 | 0-1011-1-1    | .1111....1....1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   704 | 1-0111-1-1    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   705 | 11-111-1-1    | .........1..............1....... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   706 | 10-0000--1    | ...11........................... 1 . . . ...  . . . .  . 1. .1 .1 .1 1 1  . . . .......... ... .      |
--   707 | 0--1000--1    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . ...1....1. ... .      |
--   708 | 10-0100--1    | ................................ . . . . ...  . 1 . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   709 | -1-1100--1    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   710 | -1-0010--1    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   711 | 10-00-0--1    | ..1............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   712 | -1111-0--1    | ................................ . . . . ...  1 1 . 1  . .. .. .. .. . .  . . . .......... ... .      |
--   713 | 01-1011--1    | .11111....1...........1..1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   714 | 1-1-011--1    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   715 | 11-1111--1    | ................................ . . . . ...  . 1 1 1  . .1 .. .. .. . 1  . . . .......... ... .      |
--   716 | -11-111--1    | 1...11.........1..........1...1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   717 | 011-1-1--1    | .1111.....1............1..1..... . . . . ...  . . . .  . .. .1 .1 .. . .  1 . . .......... ... .      |
--   718 | 1-10--1--1    | ................................ 1 . . . ...  . . 1 .  1 .1 .1 .. .1 1 1  . . . .......... ... .      |
--   719 | 10-010---1    | 1............................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   720 | 10-001---1    | 1............................... . . . . ...  . 1 . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   721 | 1-10-----1    | 1..111....1.........1.....1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   722 | 0-1100000-    | .1.1.1....................11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   723 | 01-100000-    | ..111.....1.......11..11..11..11 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   724 | 010010000-    | ..111.....1.......11..11..11..11 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   725 | 000110000-    | ................................ . . . . ...  . 1 1 .  . .. .. .. .. . .  . 1 . ...1.1.11. ... .      |
--   726 | 01-110000-    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   727 | -010-0000-    | ................................ . . . . ...  1 . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   728 | 010001000-    | ..111.....1.........1111....1111 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   729 | 11011-000-    | ................................ . . . . ...  . . . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   730 | 1--11-000-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   731 | 011-1-000-    | .1.1.1.........1.............11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   732 | 11-0--000-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . 11.....1.. ... .      |
--   733 | 0-0000100-    | ..111.....1.......11..11..11..11 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   734 | -0-000100-    | ................................ . . . . ...  . . . .  . .. .1 .. .1 1 .  . . . .......... ... .      |
--   735 | 01-100100-    | ..111.....1.........1111....1111 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   736 | 1-1-00100-    | 1..111....1........1....11111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   737 | --1-00100-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   738 | 010010100-    | ..111.....1.........1111....1111 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   739 | 0-1101100-    | ..........1...1..........1..1... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   740 | 01-101100-    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   741 | 100-11100-    | .11.1....1...................... 1 . . . ...  . 1 . .  . .. 1. .. .. . .  . . . .......... ... .      |
--   742 | 1--0-1100-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   743 | -011-1100-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . 1.1111.1.1 ... .      |
--   744 | -0100-100-    | .1.1..........1.1...........111. . . . . ...  1 . 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   745 | -01000-00-    | ................................ . . . . ...  . . 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   746 | 11-000-00-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   747 | 000001-00-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   748 | 0-1011-00-    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . ..1.1.111. ... .      |
--   749 | 0--111-00-    | ................................ . . . . ...  . 1 . 1  . .. .. .. .. . .  . . . .......... ... .      |
--   750 | 110-11-00-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . ....1.1.1. ... .      |
--   751 | --1-11-00-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   752 | ---0---00-    | ................................ . . . . 1.1  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   753 | 0-1100010-    | .1...1...1....1.........11.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   754 | 00-010010-    | ................................ . . . . ...  . . 1 .  . .. .. .. .. . .  . 1 . ..1.1...1. ... .      |
--   755 | 0000-0010-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   756 | 11-001010-    | ................................ . . . . ...  1 . 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   757 | -1-1-1010-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   758 | -1111-010-    | ................................ . . . . ...  . 1 1 1  . .. .. .. .. . .  . . . .......... ... .      |
--   759 | 101---010-    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   760 | 1--000110-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   761 | 110100110-    | .1.1.1....1...1...........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   762 | -00-10110-    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . ....1...1. ... .      |
--   763 | 01---0110-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   764 | 0--001110-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . ..1..11.11 ... .      |
--   765 | 00011-110-    | ................................ . . . . ...  . . 1 .  . .. .. .. .. . .  . 1 . ...1...... ... .      |
--   766 | 10011-110-    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   767 | 10-100-10-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . ...1..1... ... .      |
--   768 | ----01-10-    | ................................ . . . . 1.1  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   769 | 000111-10-    | .1.1.1........1.1...........111. . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   770 | 11-111-10-    | 1...11....1........11...1.111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   771 | 01-0-1-10-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   772 | -1-0-00-0-    | ................................ . . . . ...  . . 1 .  . .. .. .. .. . .  . . . .....1...1 ... .      |
--   773 | -110110-0-    | ................................ . . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   774 | 01-1-10-0-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   775 | 0-0-1-0-0-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   776 | -010001-0-    | .1.1..........1.1...........111. . . . . ...  1 . 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   777 | 1101001-0-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . 11.1...11. ... .      |
--   778 | 10-10-1-0-    | ................................ . . . . ...  . 1 1 1  . .. .. .. .. . .  . . 1 1........1 ... .      |
--   779 | --0111--0-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   780 | 0-111---0-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   781 | -01000001-    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   782 | 110100001-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   783 | -01010001-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . 1 . .......... 1.1 .      |
--   784 | 11-010001-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . 11..1....1 ... .      |
--   785 | 10--10001-    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   786 | 0-00-0001-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   787 | -0-1-0001-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   788 | -0-001001-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   789 | -0--01001-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   790 | 000-11001-    | ................................ 1 . . . ...  . . . .  . 1. .1 .1 .1 1 1  . . . .......... ... .      |
--   791 | -1--11001-    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   792 | 0001-1001-    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   793 | -1-11-001-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   794 | -00100101-    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   795 | 0001-0101-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . 1 . .......... 1.. .      |
--   796 | 00-011101-    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   797 | 100-11101-    | ..111....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   798 | 1-1-0-101-    | 1..111...................11111.. . . . . ...  1 . . 1  . .. 1. 11 .. . .  . . . .......... ... .      |
--   799 | -1--0-101-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   800 | --1-1-101-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   801 | -00001-01-    | .11.1........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   802 | 0-0001-01-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   803 | ---111-01-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   804 | 000100011-    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   805 | 01-110011-    | ..............1................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   806 | 0000-0011-    | ................................ . . . . ...  . 1 . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   807 | -000-0011-    | ................................ . 1 . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   808 | 0-00-0011-    | .11.1........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   809 | 10-1-0011-    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   810 | -0-1-0011-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... 1.. .      |
--   811 | 01-101011-    | .11111..............1.....111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   812 | 0000-1011-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   813 | 0100-1011-    | .11111.............1......111... 1 . . . ...  . . 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   814 | -1-01-011-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   815 | -1--1-011-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   816 | 1---00111-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   817 | 00-010111-    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . 1 . .......... 1.1 .      |
--   818 | ---110111-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   819 | 11--10111-    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   820 | 1101-0111-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   821 | 000101111-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . 1 . .......... 1.. .      |
--   822 | 01-101111-    | .1111................111111..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   823 | --1-11111-    | .....1........1....11....1.1.... 1 . . . ...  . 1 1 .  . 1. .. .. .. . 1  . . . .......... ... .      |
--   824 | -11--1111-    | .11111....1........1..11.1111... 1 . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   825 | --1--1111-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   826 | -111--111-    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   827 | 101--0-11-    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   828 | 01-101-11-    | ................................ 1 . . . ...  . 1 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   829 | 1-1-01-11-    | ................................ . . . . ...  . . . .  . .. 1. 11 .. . .  . . . .......... ... .      |
--   830 | --1-11-11-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   831 | ---0-1-11-    | ................................ . . . . ..1  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   832 | -111-1-11-    | 1...11.........1.........11111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   833 | 1--1-1-11-    | ................................ . . . . ...  1 . . 1  . .. .. .. .. . .  . . . .1....1... ... .      |
--   834 | 1-1-000-1-    | 1..111.........1..........11..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   835 | 10-0110-1-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   836 | 1-01-10-1-    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . ...1.....1 ... .      |
--   837 | 1-0-101-1-    | ................................ . . . . ...  1 1 . 1  . .. .. .. .. . .  . . . 11.11.1..1 1.. .      |
--   838 | 111-101-1-    | ................................ . . . . ...  1 1 . 1  . .. .. .1 .. . .  . . . .......... ... .      |
--   839 | -----01-1-    | ................................ . . . . .11  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   840 | -000011-1-    | ................................ . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   841 | 11-1111-1-    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   842 | 101--11-1-    | ................................ . . . . ...  . 1 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   843 | 01---11-1-    | ................................ . . . . ...  . 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   844 | 10-00-1-1-    | ................................ 1 . . . ...  . 1 . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   845 | -1101-1-1-    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   846 | 011-1-1-1-    | .11111...1.....1......111.1..11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   847 | -00010--1-    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   848 | -011-0--1-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   849 | 10-001--1-    | .11.1........................... 1 . . . ...  . 1 . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   850 | -1--11--1-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   851 | 0100----1-    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   852 | 10-01000--    | .11.1........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   853 | -110-000--    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   854 | 00011100--    | .11111.........1......1....1.1.. 1 . . . ...  . . 1 .  . 1. .. .. .. . .  . . . .......... ... .      |
--   855 | 00000010--    | .11111....................111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   856 | -0100010--    | .1.1.1........1...........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   857 | 00-00010--    | ................................ . . . . ...  1 . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   858 | --101110--    | 1..111....1...............1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   859 | 1101-110--    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . .1.1..1... 1.1 .      |
--   860 | 0-001-10--    | ................................ . . . . ...  1 . 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   861 | 100110-0--    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . 1....11111 ... .      |
--   862 | -1--11-0--    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   863 | 01-----0--    | ................................ . . . . ...  1 . 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   864 | -0100101--    | .1.1.1........1...........11111. . . . . ...  1 . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   865 | -1100101--    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   866 | 100-1101--    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . 1...11..1. ... .      |
--   867 | 11011-01--    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . 11.11..1.. 1.1 .      |
--   868 | ---01011--    | ................................ . . . . ...  1 . 1 .  . .. .. .. .. . .  . . . ......1... ... .      |
--   869 | --110111--    | .1111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   870 | -0011111--    | .1.1.1........1.11........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   871 | -100-111--    | ................................ . . . . ...  1 1 . 1  . .. .. .. .. . .  . . . .......... ... .      |
--   872 | 1-1--111--    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   873 | -1101-11--    | 1...11....1...............1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   874 | -1-11-11--    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   875 | 0--11-11--    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   876 | ----10-1--    | ................................ . . . . 1..  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   877 | 0100-0-1--    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   878 | --0111-1--    | ................................ . . . . ...  1 . . .  . .. .. .. .. . .  . . . ...1...... ... .      |
--   879 | ---11--1--    | ................................ . . . . .1.  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   880 | 0-11-10---    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   881 | ----0-0---    | ................................ . . . . 1..  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   882 | ----111---    | ................................ . . . . 11.  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   883 | 11011-1---    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   884 | ----00----    | ................................ . . . . .1.  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   885 | ---111----    | ................................ . . . . .1.  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   886 | 111-------    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   887 | --1-------    | ................................ . . . . 1.1  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   888 | -1--------    | ................................ . . . . 111  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   889 | 0---------    | ................................ . . . . 111  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   890 | ----------    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... .1. .      |
--      *=======================================================================================================================*
--
-- Table ROM64_INSTR Signal Assignments for Product Terms
MQQ1:ROM64_INSTR_PT(1) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100000000"));
MQQ2:ROM64_INSTR_PT(2) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000000"));
MQQ3:ROM64_INSTR_PT(3) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000000"));
MQQ4:ROM64_INSTR_PT(4) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000000"));
MQQ5:ROM64_INSTR_PT(5) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000000"));
MQQ6:ROM64_INSTR_PT(6) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110000000"));
MQQ7:ROM64_INSTR_PT(7) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000000"));
MQQ8:ROM64_INSTR_PT(8) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00100000"));
MQQ9:ROM64_INSTR_PT(9) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100000"));
MQQ10:ROM64_INSTR_PT(10) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100000"));
MQQ11:ROM64_INSTR_PT(11) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100000"));
MQQ12:ROM64_INSTR_PT(12) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000000"));
MQQ13:ROM64_INSTR_PT(13) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000000"));
MQQ14:ROM64_INSTR_PT(14) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010000"));
MQQ15:ROM64_INSTR_PT(15) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010000"));
MQQ16:ROM64_INSTR_PT(16) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101010000"));
MQQ17:ROM64_INSTR_PT(17) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000110000"));
MQQ18:ROM64_INSTR_PT(18) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010110000"));
MQQ19:ROM64_INSTR_PT(19) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0110000"));
MQQ20:ROM64_INSTR_PT(20) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110000"));
MQQ21:ROM64_INSTR_PT(21) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110000"));
MQQ22:ROM64_INSTR_PT(22) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110000"));
MQQ23:ROM64_INSTR_PT(23) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010000"));
MQQ24:ROM64_INSTR_PT(24) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110000"));
MQQ25:ROM64_INSTR_PT(25) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ26:ROM64_INSTR_PT(26) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000000"));
MQQ27:ROM64_INSTR_PT(27) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100000"));
MQQ28:ROM64_INSTR_PT(28) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010000"));
MQQ29:ROM64_INSTR_PT(29) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110000"));
MQQ30:ROM64_INSTR_PT(30) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ31:ROM64_INSTR_PT(31) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110000"));
MQQ32:ROM64_INSTR_PT(32) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0010000"));
MQQ33:ROM64_INSTR_PT(33) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010000"));
MQQ34:ROM64_INSTR_PT(34) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010000"));
MQQ35:ROM64_INSTR_PT(35) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110000"));
MQQ36:ROM64_INSTR_PT(36) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001000"));
MQQ37:ROM64_INSTR_PT(37) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101001000"));
MQQ38:ROM64_INSTR_PT(38) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110001000"));
MQQ39:ROM64_INSTR_PT(39) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001000"));
MQQ40:ROM64_INSTR_PT(40) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101000"));
MQQ41:ROM64_INSTR_PT(41) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001101000"));
MQQ42:ROM64_INSTR_PT(42) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101000"));
MQQ43:ROM64_INSTR_PT(43) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101000"));
MQQ44:ROM64_INSTR_PT(44) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101000"));
MQQ45:ROM64_INSTR_PT(45) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111101000"));
MQQ46:ROM64_INSTR_PT(46) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001000"));
MQQ47:ROM64_INSTR_PT(47) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101000"));
MQQ48:ROM64_INSTR_PT(48) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001011000"));
MQQ49:ROM64_INSTR_PT(49) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011011000"));
MQQ50:ROM64_INSTR_PT(50) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011000"));
MQQ51:ROM64_INSTR_PT(51) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111000"));
MQQ52:ROM64_INSTR_PT(52) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111000"));
MQQ53:ROM64_INSTR_PT(53) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111000"));
MQQ54:ROM64_INSTR_PT(54) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011000"));
MQQ55:ROM64_INSTR_PT(55) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111000"));
MQQ56:ROM64_INSTR_PT(56) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111000"));
MQQ57:ROM64_INSTR_PT(57) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111000"));
MQQ58:ROM64_INSTR_PT(58) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001000"));
MQQ59:ROM64_INSTR_PT(59) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011000"));
MQQ60:ROM64_INSTR_PT(60) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011000"));
MQQ61:ROM64_INSTR_PT(61) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100111000"));
MQQ62:ROM64_INSTR_PT(62) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111000"));
MQQ63:ROM64_INSTR_PT(63) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000000"));
MQQ64:ROM64_INSTR_PT(64) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000000"));
MQQ65:ROM64_INSTR_PT(65) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000000"));
MQQ66:ROM64_INSTR_PT(66) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010000"));
MQQ67:ROM64_INSTR_PT(67) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ68:ROM64_INSTR_PT(68) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100000"));
MQQ69:ROM64_INSTR_PT(69) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010000"));
MQQ70:ROM64_INSTR_PT(70) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001000"));
MQQ71:ROM64_INSTR_PT(71) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011000"));
MQQ72:ROM64_INSTR_PT(72) <=
    Eq(( ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000"));
MQQ73:ROM64_INSTR_PT(73) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100000100"));
MQQ74:ROM64_INSTR_PT(74) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000100"));
MQQ75:ROM64_INSTR_PT(75) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000100"));
MQQ76:ROM64_INSTR_PT(76) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000100"));
MQQ77:ROM64_INSTR_PT(77) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000100"));
MQQ78:ROM64_INSTR_PT(78) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000100"));
MQQ79:ROM64_INSTR_PT(79) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000100"));
MQQ80:ROM64_INSTR_PT(80) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100100100"));
MQQ81:ROM64_INSTR_PT(81) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100100"));
MQQ82:ROM64_INSTR_PT(82) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100100"));
MQQ83:ROM64_INSTR_PT(83) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100100"));
MQQ84:ROM64_INSTR_PT(84) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11100100"));
MQQ85:ROM64_INSTR_PT(85) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100100"));
MQQ86:ROM64_INSTR_PT(86) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000100"));
MQQ87:ROM64_INSTR_PT(87) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000100"));
MQQ88:ROM64_INSTR_PT(88) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100100"));
MQQ89:ROM64_INSTR_PT(89) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100010100"));
MQQ90:ROM64_INSTR_PT(90) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110010100"));
MQQ91:ROM64_INSTR_PT(91) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010100"));
MQQ92:ROM64_INSTR_PT(92) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010100"));
MQQ93:ROM64_INSTR_PT(93) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010100"));
MQQ94:ROM64_INSTR_PT(94) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010100"));
MQQ95:ROM64_INSTR_PT(95) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000110100"));
MQQ96:ROM64_INSTR_PT(96) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010110100"));
MQQ97:ROM64_INSTR_PT(97) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110100"));
MQQ98:ROM64_INSTR_PT(98) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110100"));
MQQ99:ROM64_INSTR_PT(99) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110100"));
MQQ100:ROM64_INSTR_PT(100) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110100"));
MQQ101:ROM64_INSTR_PT(101) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110100"));
MQQ102:ROM64_INSTR_PT(102) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000100"));
MQQ103:ROM64_INSTR_PT(103) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010100"));
MQQ104:ROM64_INSTR_PT(104) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110100"));
MQQ105:ROM64_INSTR_PT(105) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010100"));
MQQ106:ROM64_INSTR_PT(106) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100001100"));
MQQ107:ROM64_INSTR_PT(107) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001001100"));
MQQ108:ROM64_INSTR_PT(108) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001001100"));
MQQ109:ROM64_INSTR_PT(109) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001100"));
MQQ110:ROM64_INSTR_PT(110) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001100"));
MQQ111:ROM64_INSTR_PT(111) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001100"));
MQQ112:ROM64_INSTR_PT(112) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101100"));
MQQ113:ROM64_INSTR_PT(113) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100101100"));
MQQ114:ROM64_INSTR_PT(114) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010101100"));
MQQ115:ROM64_INSTR_PT(115) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101100"));
MQQ116:ROM64_INSTR_PT(116) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101100"));
MQQ117:ROM64_INSTR_PT(117) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ118:ROM64_INSTR_PT(118) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ119:ROM64_INSTR_PT(119) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011100"));
MQQ120:ROM64_INSTR_PT(120) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011100"));
MQQ121:ROM64_INSTR_PT(121) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011011100"));
MQQ122:ROM64_INSTR_PT(122) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ123:ROM64_INSTR_PT(123) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100111100"));
MQQ124:ROM64_INSTR_PT(124) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111100"));
MQQ125:ROM64_INSTR_PT(125) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ126:ROM64_INSTR_PT(126) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ127:ROM64_INSTR_PT(127) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011100"));
MQQ128:ROM64_INSTR_PT(128) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011100"));
MQQ129:ROM64_INSTR_PT(129) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111100"));
MQQ130:ROM64_INSTR_PT(130) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ131:ROM64_INSTR_PT(131) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011100"));
MQQ132:ROM64_INSTR_PT(132) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ133:ROM64_INSTR_PT(133) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001100"));
MQQ134:ROM64_INSTR_PT(134) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101100"));
MQQ135:ROM64_INSTR_PT(135) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ136:ROM64_INSTR_PT(136) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111100"));
MQQ137:ROM64_INSTR_PT(137) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111100"));
MQQ138:ROM64_INSTR_PT(138) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0100100"));
MQQ139:ROM64_INSTR_PT(139) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010100"));
MQQ140:ROM64_INSTR_PT(140) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010100"));
MQQ141:ROM64_INSTR_PT(141) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001100"));
MQQ142:ROM64_INSTR_PT(142) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001100"));
MQQ143:ROM64_INSTR_PT(143) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ144:ROM64_INSTR_PT(144) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111100"));
MQQ145:ROM64_INSTR_PT(145) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ146:ROM64_INSTR_PT(146) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001100"));
MQQ147:ROM64_INSTR_PT(147) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000000"));
MQQ148:ROM64_INSTR_PT(148) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010000"));
MQQ149:ROM64_INSTR_PT(149) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010000"));
MQQ150:ROM64_INSTR_PT(150) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001000"));
MQQ151:ROM64_INSTR_PT(151) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001000"));
MQQ152:ROM64_INSTR_PT(152) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1000"));
MQQ153:ROM64_INSTR_PT(153) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000100"));
MQQ154:ROM64_INSTR_PT(154) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000100"));
MQQ155:ROM64_INSTR_PT(155) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100100"));
MQQ156:ROM64_INSTR_PT(156) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("00100"));
MQQ157:ROM64_INSTR_PT(157) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ158:ROM64_INSTR_PT(158) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ159:ROM64_INSTR_PT(159) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111100"));
MQQ160:ROM64_INSTR_PT(160) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011100"));
MQQ161:ROM64_INSTR_PT(161) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011100"));
MQQ162:ROM64_INSTR_PT(162) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111100"));
MQQ163:ROM64_INSTR_PT(163) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("01000"));
MQQ164:ROM64_INSTR_PT(164) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000100"));
MQQ165:ROM64_INSTR_PT(165) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("10100"));
MQQ166:ROM64_INSTR_PT(166) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ167:ROM64_INSTR_PT(167) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("01100"));
MQQ168:ROM64_INSTR_PT(168) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100000010"));
MQQ169:ROM64_INSTR_PT(169) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000010"));
MQQ170:ROM64_INSTR_PT(170) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000010"));
MQQ171:ROM64_INSTR_PT(171) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000010"));
MQQ172:ROM64_INSTR_PT(172) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000010"));
MQQ173:ROM64_INSTR_PT(173) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100010"));
MQQ174:ROM64_INSTR_PT(174) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100010"));
MQQ175:ROM64_INSTR_PT(175) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100010"));
MQQ176:ROM64_INSTR_PT(176) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000010"));
MQQ177:ROM64_INSTR_PT(177) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ178:ROM64_INSTR_PT(178) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("000010"));
MQQ179:ROM64_INSTR_PT(179) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010010"));
MQQ180:ROM64_INSTR_PT(180) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001110010"));
MQQ181:ROM64_INSTR_PT(181) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110010"));
MQQ182:ROM64_INSTR_PT(182) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110010"));
MQQ183:ROM64_INSTR_PT(183) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110010"));
MQQ184:ROM64_INSTR_PT(184) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010010"));
MQQ185:ROM64_INSTR_PT(185) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010010"));
MQQ186:ROM64_INSTR_PT(186) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110010"));
MQQ187:ROM64_INSTR_PT(187) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110010"));
MQQ188:ROM64_INSTR_PT(188) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ189:ROM64_INSTR_PT(189) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000010"));
MQQ190:ROM64_INSTR_PT(190) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000010"));
MQQ191:ROM64_INSTR_PT(191) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100010"));
MQQ192:ROM64_INSTR_PT(192) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ193:ROM64_INSTR_PT(193) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110010"));
MQQ194:ROM64_INSTR_PT(194) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110010"));
MQQ195:ROM64_INSTR_PT(195) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110010"));
MQQ196:ROM64_INSTR_PT(196) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ197:ROM64_INSTR_PT(197) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110010"));
MQQ198:ROM64_INSTR_PT(198) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ199:ROM64_INSTR_PT(199) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001010"));
MQQ200:ROM64_INSTR_PT(200) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101001010"));
MQQ201:ROM64_INSTR_PT(201) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001001010"));
MQQ202:ROM64_INSTR_PT(202) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001010"));
MQQ203:ROM64_INSTR_PT(203) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001010"));
MQQ204:ROM64_INSTR_PT(204) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001010"));
MQQ205:ROM64_INSTR_PT(205) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101010"));
MQQ206:ROM64_INSTR_PT(206) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101010"));
MQQ207:ROM64_INSTR_PT(207) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101010"));
MQQ208:ROM64_INSTR_PT(208) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101010"));
MQQ209:ROM64_INSTR_PT(209) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101010"));
MQQ210:ROM64_INSTR_PT(210) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001010"));
MQQ211:ROM64_INSTR_PT(211) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011010"));
MQQ212:ROM64_INSTR_PT(212) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ213:ROM64_INSTR_PT(213) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011010"));
MQQ214:ROM64_INSTR_PT(214) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011011010"));
MQQ215:ROM64_INSTR_PT(215) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111010"));
MQQ216:ROM64_INSTR_PT(216) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011111010"));
MQQ217:ROM64_INSTR_PT(217) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111010"));
MQQ218:ROM64_INSTR_PT(218) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111010"));
MQQ219:ROM64_INSTR_PT(219) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011010"));
MQQ220:ROM64_INSTR_PT(220) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011010"));
MQQ221:ROM64_INSTR_PT(221) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100111010"));
MQQ222:ROM64_INSTR_PT(222) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111010"));
MQQ223:ROM64_INSTR_PT(223) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111010"));
MQQ224:ROM64_INSTR_PT(224) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101010"));
MQQ225:ROM64_INSTR_PT(225) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011010"));
MQQ226:ROM64_INSTR_PT(226) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ227:ROM64_INSTR_PT(227) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011010"));
MQQ228:ROM64_INSTR_PT(228) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100010"));
MQQ229:ROM64_INSTR_PT(229) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100010"));
MQQ230:ROM64_INSTR_PT(230) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010010"));
MQQ231:ROM64_INSTR_PT(231) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ232:ROM64_INSTR_PT(232) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001010"));
MQQ233:ROM64_INSTR_PT(233) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101010"));
MQQ234:ROM64_INSTR_PT(234) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011010"));
MQQ235:ROM64_INSTR_PT(235) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011010"));
MQQ236:ROM64_INSTR_PT(236) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100000110"));
MQQ237:ROM64_INSTR_PT(237) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110000110"));
MQQ238:ROM64_INSTR_PT(238) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000110"));
MQQ239:ROM64_INSTR_PT(239) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000110"));
MQQ240:ROM64_INSTR_PT(240) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000110"));
MQQ241:ROM64_INSTR_PT(241) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000110"));
MQQ242:ROM64_INSTR_PT(242) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111000110"));
MQQ243:ROM64_INSTR_PT(243) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000110"));
MQQ244:ROM64_INSTR_PT(244) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000110"));
MQQ245:ROM64_INSTR_PT(245) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000100110"));
MQQ246:ROM64_INSTR_PT(246) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100110"));
MQQ247:ROM64_INSTR_PT(247) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001100110"));
MQQ248:ROM64_INSTR_PT(248) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000110"));
MQQ249:ROM64_INSTR_PT(249) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000110"));
MQQ250:ROM64_INSTR_PT(250) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000110"));
MQQ251:ROM64_INSTR_PT(251) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100110"));
MQQ252:ROM64_INSTR_PT(252) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110010110"));
MQQ253:ROM64_INSTR_PT(253) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010110"));
MQQ254:ROM64_INSTR_PT(254) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010110"));
MQQ255:ROM64_INSTR_PT(255) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110110"));
MQQ256:ROM64_INSTR_PT(256) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110110"));
MQQ257:ROM64_INSTR_PT(257) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110110"));
MQQ258:ROM64_INSTR_PT(258) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110110"));
MQQ259:ROM64_INSTR_PT(259) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100110110"));
MQQ260:ROM64_INSTR_PT(260) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110110"));
MQQ261:ROM64_INSTR_PT(261) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110110"));
MQQ262:ROM64_INSTR_PT(262) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100110"));
MQQ263:ROM64_INSTR_PT(263) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100110110"));
MQQ264:ROM64_INSTR_PT(264) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110110"));
MQQ265:ROM64_INSTR_PT(265) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100001110"));
MQQ266:ROM64_INSTR_PT(266) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001110"));
MQQ267:ROM64_INSTR_PT(267) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110001110"));
MQQ268:ROM64_INSTR_PT(268) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001110"));
MQQ269:ROM64_INSTR_PT(269) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001110"));
MQQ270:ROM64_INSTR_PT(270) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000101110"));
MQQ271:ROM64_INSTR_PT(271) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100101110"));
MQQ272:ROM64_INSTR_PT(272) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101110"));
MQQ273:ROM64_INSTR_PT(273) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101110"));
MQQ274:ROM64_INSTR_PT(274) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101110"));
MQQ275:ROM64_INSTR_PT(275) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101110"));
MQQ276:ROM64_INSTR_PT(276) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101110"));
MQQ277:ROM64_INSTR_PT(277) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011110"));
MQQ278:ROM64_INSTR_PT(278) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011110"));
MQQ279:ROM64_INSTR_PT(279) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ280:ROM64_INSTR_PT(280) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111110"));
MQQ281:ROM64_INSTR_PT(281) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111110"));
MQQ282:ROM64_INSTR_PT(282) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111110"));
MQQ283:ROM64_INSTR_PT(283) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011110"));
MQQ284:ROM64_INSTR_PT(284) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011110"));
MQQ285:ROM64_INSTR_PT(285) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ286:ROM64_INSTR_PT(286) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111110"));
MQQ287:ROM64_INSTR_PT(287) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111110"));
MQQ288:ROM64_INSTR_PT(288) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111110"));
MQQ289:ROM64_INSTR_PT(289) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111110"));
MQQ290:ROM64_INSTR_PT(290) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ291:ROM64_INSTR_PT(291) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111110"));
MQQ292:ROM64_INSTR_PT(292) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111110"));
MQQ293:ROM64_INSTR_PT(293) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ294:ROM64_INSTR_PT(294) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110110"));
MQQ295:ROM64_INSTR_PT(295) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100110"));
MQQ296:ROM64_INSTR_PT(296) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001110"));
MQQ297:ROM64_INSTR_PT(297) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ298:ROM64_INSTR_PT(298) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111110"));
MQQ299:ROM64_INSTR_PT(299) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011110"));
MQQ300:ROM64_INSTR_PT(300) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ301:ROM64_INSTR_PT(301) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101110"));
MQQ302:ROM64_INSTR_PT(302) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101110"));
MQQ303:ROM64_INSTR_PT(303) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000010"));
MQQ304:ROM64_INSTR_PT(304) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011010"));
MQQ305:ROM64_INSTR_PT(305) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ306:ROM64_INSTR_PT(306) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ307:ROM64_INSTR_PT(307) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101010"));
MQQ308:ROM64_INSTR_PT(308) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000110"));
MQQ309:ROM64_INSTR_PT(309) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000110"));
MQQ310:ROM64_INSTR_PT(310) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010110"));
MQQ311:ROM64_INSTR_PT(311) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110110"));
MQQ312:ROM64_INSTR_PT(312) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001110"));
MQQ313:ROM64_INSTR_PT(313) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001110"));
MQQ314:ROM64_INSTR_PT(314) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111110"));
MQQ315:ROM64_INSTR_PT(315) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ316:ROM64_INSTR_PT(316) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010110"));
MQQ317:ROM64_INSTR_PT(317) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010010"));
MQQ318:ROM64_INSTR_PT(318) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("01010"));
MQQ319:ROM64_INSTR_PT(319) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ320:ROM64_INSTR_PT(320) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0000010"));
MQQ321:ROM64_INSTR_PT(321) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000000"));
MQQ322:ROM64_INSTR_PT(322) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010000"));
MQQ323:ROM64_INSTR_PT(323) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000000"));
MQQ324:ROM64_INSTR_PT(324) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101000"));
MQQ325:ROM64_INSTR_PT(325) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101000"));
MQQ326:ROM64_INSTR_PT(326) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101000"));
MQQ327:ROM64_INSTR_PT(327) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100000"));
MQQ328:ROM64_INSTR_PT(328) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011000"));
MQQ329:ROM64_INSTR_PT(329) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0000100"));
MQQ330:ROM64_INSTR_PT(330) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000100"));
MQQ331:ROM64_INSTR_PT(331) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000100"));
MQQ332:ROM64_INSTR_PT(332) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000100"));
MQQ333:ROM64_INSTR_PT(333) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001100"));
MQQ334:ROM64_INSTR_PT(334) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00101100"));
MQQ335:ROM64_INSTR_PT(335) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011100"));
MQQ336:ROM64_INSTR_PT(336) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000000"));
MQQ337:ROM64_INSTR_PT(337) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ338:ROM64_INSTR_PT(338) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000010"));
MQQ339:ROM64_INSTR_PT(339) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ340:ROM64_INSTR_PT(340) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010010"));
MQQ341:ROM64_INSTR_PT(341) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ342:ROM64_INSTR_PT(342) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ343:ROM64_INSTR_PT(343) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001010"));
MQQ344:ROM64_INSTR_PT(344) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001010"));
MQQ345:ROM64_INSTR_PT(345) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100110"));
MQQ346:ROM64_INSTR_PT(346) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ347:ROM64_INSTR_PT(347) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ348:ROM64_INSTR_PT(348) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ349:ROM64_INSTR_PT(349) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101110"));
MQQ350:ROM64_INSTR_PT(350) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ351:ROM64_INSTR_PT(351) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101010"));
MQQ352:ROM64_INSTR_PT(352) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101110"));
MQQ353:ROM64_INSTR_PT(353) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011110"));
MQQ354:ROM64_INSTR_PT(354) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000000"));
MQQ355:ROM64_INSTR_PT(355) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ356:ROM64_INSTR_PT(356) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000010"));
MQQ357:ROM64_INSTR_PT(357) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100010"));
MQQ358:ROM64_INSTR_PT(358) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110110"));
MQQ359:ROM64_INSTR_PT(359) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011110"));
MQQ360:ROM64_INSTR_PT(360) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100010"));
MQQ361:ROM64_INSTR_PT(361) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100000001"));
MQQ362:ROM64_INSTR_PT(362) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000001"));
MQQ363:ROM64_INSTR_PT(363) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000001"));
MQQ364:ROM64_INSTR_PT(364) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110000001"));
MQQ365:ROM64_INSTR_PT(365) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000001"));
MQQ366:ROM64_INSTR_PT(366) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100001"));
MQQ367:ROM64_INSTR_PT(367) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11100001"));
MQQ368:ROM64_INSTR_PT(368) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000001"));
MQQ369:ROM64_INSTR_PT(369) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ370:ROM64_INSTR_PT(370) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010001"));
MQQ371:ROM64_INSTR_PT(371) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010001"));
MQQ372:ROM64_INSTR_PT(372) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010001"));
MQQ373:ROM64_INSTR_PT(373) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110001"));
MQQ374:ROM64_INSTR_PT(374) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010110001"));
MQQ375:ROM64_INSTR_PT(375) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001110001"));
MQQ376:ROM64_INSTR_PT(376) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00110001"));
MQQ377:ROM64_INSTR_PT(377) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110001"));
MQQ378:ROM64_INSTR_PT(378) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110001"));
MQQ379:ROM64_INSTR_PT(379) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110001"));
MQQ380:ROM64_INSTR_PT(380) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110001"));
MQQ381:ROM64_INSTR_PT(381) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110001"));
MQQ382:ROM64_INSTR_PT(382) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110001"));
MQQ383:ROM64_INSTR_PT(383) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ384:ROM64_INSTR_PT(384) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100001"));
MQQ385:ROM64_INSTR_PT(385) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100110001"));
MQQ386:ROM64_INSTR_PT(386) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110001"));
MQQ387:ROM64_INSTR_PT(387) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010001"));
MQQ388:ROM64_INSTR_PT(388) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001001"));
MQQ389:ROM64_INSTR_PT(389) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111001001"));
MQQ390:ROM64_INSTR_PT(390) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001001"));
MQQ391:ROM64_INSTR_PT(391) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001001"));
MQQ392:ROM64_INSTR_PT(392) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101001"));
MQQ393:ROM64_INSTR_PT(393) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00101001"));
MQQ394:ROM64_INSTR_PT(394) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101001"));
MQQ395:ROM64_INSTR_PT(395) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001101001"));
MQQ396:ROM64_INSTR_PT(396) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101001"));
MQQ397:ROM64_INSTR_PT(397) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101001"));
MQQ398:ROM64_INSTR_PT(398) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111101001"));
MQQ399:ROM64_INSTR_PT(399) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001001"));
MQQ400:ROM64_INSTR_PT(400) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("001001"));
MQQ401:ROM64_INSTR_PT(401) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011001"));
MQQ402:ROM64_INSTR_PT(402) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001011001"));
MQQ403:ROM64_INSTR_PT(403) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011111001"));
MQQ404:ROM64_INSTR_PT(404) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111001"));
MQQ405:ROM64_INSTR_PT(405) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011001"));
MQQ406:ROM64_INSTR_PT(406) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011001"));
MQQ407:ROM64_INSTR_PT(407) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011001"));
MQQ408:ROM64_INSTR_PT(408) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111001"));
MQQ409:ROM64_INSTR_PT(409) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111001"));
MQQ410:ROM64_INSTR_PT(410) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111001"));
MQQ411:ROM64_INSTR_PT(411) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011001"));
MQQ412:ROM64_INSTR_PT(412) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111001"));
MQQ413:ROM64_INSTR_PT(413) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111001"));
MQQ414:ROM64_INSTR_PT(414) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000001"));
MQQ415:ROM64_INSTR_PT(415) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ416:ROM64_INSTR_PT(416) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100001"));
MQQ417:ROM64_INSTR_PT(417) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010001"));
MQQ418:ROM64_INSTR_PT(418) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010001"));
MQQ419:ROM64_INSTR_PT(419) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101001"));
MQQ420:ROM64_INSTR_PT(420) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011001"));
MQQ421:ROM64_INSTR_PT(421) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011001"));
MQQ422:ROM64_INSTR_PT(422) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100000101"));
MQQ423:ROM64_INSTR_PT(423) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000101"));
MQQ424:ROM64_INSTR_PT(424) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000101"));
MQQ425:ROM64_INSTR_PT(425) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000101"));
MQQ426:ROM64_INSTR_PT(426) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000101"));
MQQ427:ROM64_INSTR_PT(427) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000101"));
MQQ428:ROM64_INSTR_PT(428) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000101"));
MQQ429:ROM64_INSTR_PT(429) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100100101"));
MQQ430:ROM64_INSTR_PT(430) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100101"));
MQQ431:ROM64_INSTR_PT(431) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100101"));
MQQ432:ROM64_INSTR_PT(432) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100101"));
MQQ433:ROM64_INSTR_PT(433) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100101"));
MQQ434:ROM64_INSTR_PT(434) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100101"));
MQQ435:ROM64_INSTR_PT(435) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11100101"));
MQQ436:ROM64_INSTR_PT(436) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100101"));
MQQ437:ROM64_INSTR_PT(437) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110010101"));
MQQ438:ROM64_INSTR_PT(438) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010101"));
MQQ439:ROM64_INSTR_PT(439) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101010101"));
MQQ440:ROM64_INSTR_PT(440) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010101"));
MQQ441:ROM64_INSTR_PT(441) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000110101"));
MQQ442:ROM64_INSTR_PT(442) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110101"));
MQQ443:ROM64_INSTR_PT(443) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110101"));
MQQ444:ROM64_INSTR_PT(444) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110101"));
MQQ445:ROM64_INSTR_PT(445) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110101"));
MQQ446:ROM64_INSTR_PT(446) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000101"));
MQQ447:ROM64_INSTR_PT(447) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100101"));
MQQ448:ROM64_INSTR_PT(448) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110101"));
MQQ449:ROM64_INSTR_PT(449) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110101"));
MQQ450:ROM64_INSTR_PT(450) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010101"));
MQQ451:ROM64_INSTR_PT(451) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100001101"));
MQQ452:ROM64_INSTR_PT(452) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110001101"));
MQQ453:ROM64_INSTR_PT(453) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001001101"));
MQQ454:ROM64_INSTR_PT(454) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001101"));
MQQ455:ROM64_INSTR_PT(455) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010101101"));
MQQ456:ROM64_INSTR_PT(456) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101101"));
MQQ457:ROM64_INSTR_PT(457) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101101"));
MQQ458:ROM64_INSTR_PT(458) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101101"));
MQQ459:ROM64_INSTR_PT(459) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001101"));
MQQ460:ROM64_INSTR_PT(460) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101101"));
MQQ461:ROM64_INSTR_PT(461) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011101"));
MQQ462:ROM64_INSTR_PT(462) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011101"));
MQQ463:ROM64_INSTR_PT(463) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111101"));
MQQ464:ROM64_INSTR_PT(464) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111101"));
MQQ465:ROM64_INSTR_PT(465) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011101"));
MQQ466:ROM64_INSTR_PT(466) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011101"));
MQQ467:ROM64_INSTR_PT(467) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111101"));
MQQ468:ROM64_INSTR_PT(468) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100111101"));
MQQ469:ROM64_INSTR_PT(469) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111101"));
MQQ470:ROM64_INSTR_PT(470) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111101"));
MQQ471:ROM64_INSTR_PT(471) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001101"));
MQQ472:ROM64_INSTR_PT(472) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100101"));
MQQ473:ROM64_INSTR_PT(473) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010101"));
MQQ474:ROM64_INSTR_PT(474) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110101"));
MQQ475:ROM64_INSTR_PT(475) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010101"));
MQQ476:ROM64_INSTR_PT(476) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010101"));
MQQ477:ROM64_INSTR_PT(477) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001101"));
MQQ478:ROM64_INSTR_PT(478) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001101"));
MQQ479:ROM64_INSTR_PT(479) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001101"));
MQQ480:ROM64_INSTR_PT(480) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011101"));
MQQ481:ROM64_INSTR_PT(481) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111101"));
MQQ482:ROM64_INSTR_PT(482) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ483:ROM64_INSTR_PT(483) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010001"));
MQQ484:ROM64_INSTR_PT(484) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110001"));
MQQ485:ROM64_INSTR_PT(485) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001001"));
MQQ486:ROM64_INSTR_PT(486) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001001"));
MQQ487:ROM64_INSTR_PT(487) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101001"));
MQQ488:ROM64_INSTR_PT(488) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011001"));
MQQ489:ROM64_INSTR_PT(489) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111001"));
MQQ490:ROM64_INSTR_PT(490) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111001"));
MQQ491:ROM64_INSTR_PT(491) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000101"));
MQQ492:ROM64_INSTR_PT(492) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100101"));
MQQ493:ROM64_INSTR_PT(493) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100101"));
MQQ494:ROM64_INSTR_PT(494) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100101"));
MQQ495:ROM64_INSTR_PT(495) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111101"));
MQQ496:ROM64_INSTR_PT(496) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011101"));
MQQ497:ROM64_INSTR_PT(497) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111101"));
MQQ498:ROM64_INSTR_PT(498) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101101"));
MQQ499:ROM64_INSTR_PT(499) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001101"));
MQQ500:ROM64_INSTR_PT(500) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0000001"));
MQQ501:ROM64_INSTR_PT(501) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("001101"));
MQQ502:ROM64_INSTR_PT(502) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001"));
MQQ503:ROM64_INSTR_PT(503) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100000011"));
MQQ504:ROM64_INSTR_PT(504) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000011"));
MQQ505:ROM64_INSTR_PT(505) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000011"));
MQQ506:ROM64_INSTR_PT(506) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000011"));
MQQ507:ROM64_INSTR_PT(507) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000011"));
MQQ508:ROM64_INSTR_PT(508) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010100011"));
MQQ509:ROM64_INSTR_PT(509) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100011"));
MQQ510:ROM64_INSTR_PT(510) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100011"));
MQQ511:ROM64_INSTR_PT(511) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000011"));
MQQ512:ROM64_INSTR_PT(512) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100011"));
MQQ513:ROM64_INSTR_PT(513) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000011"));
MQQ514:ROM64_INSTR_PT(514) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010011"));
MQQ515:ROM64_INSTR_PT(515) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010011"));
MQQ516:ROM64_INSTR_PT(516) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010011"));
MQQ517:ROM64_INSTR_PT(517) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010011"));
MQQ518:ROM64_INSTR_PT(518) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010011"));
MQQ519:ROM64_INSTR_PT(519) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001110011"));
MQQ520:ROM64_INSTR_PT(520) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110011"));
MQQ521:ROM64_INSTR_PT(521) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110011"));
MQQ522:ROM64_INSTR_PT(522) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110011"));
MQQ523:ROM64_INSTR_PT(523) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110011"));
MQQ524:ROM64_INSTR_PT(524) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000011"));
MQQ525:ROM64_INSTR_PT(525) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100011"));
MQQ526:ROM64_INSTR_PT(526) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100011"));
MQQ527:ROM64_INSTR_PT(527) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010011"));
MQQ528:ROM64_INSTR_PT(528) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110011"));
MQQ529:ROM64_INSTR_PT(529) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010011"));
MQQ530:ROM64_INSTR_PT(530) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001011"));
MQQ531:ROM64_INSTR_PT(531) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101001011"));
MQQ532:ROM64_INSTR_PT(532) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001001011"));
MQQ533:ROM64_INSTR_PT(533) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111001011"));
MQQ534:ROM64_INSTR_PT(534) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000101011"));
MQQ535:ROM64_INSTR_PT(535) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101011"));
MQQ536:ROM64_INSTR_PT(536) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001101011"));
MQQ537:ROM64_INSTR_PT(537) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101011"));
MQQ538:ROM64_INSTR_PT(538) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101011"));
MQQ539:ROM64_INSTR_PT(539) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001011"));
MQQ540:ROM64_INSTR_PT(540) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101011"));
MQQ541:ROM64_INSTR_PT(541) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011011"));
MQQ542:ROM64_INSTR_PT(542) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ543:ROM64_INSTR_PT(543) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011011"));
MQQ544:ROM64_INSTR_PT(544) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111011"));
MQQ545:ROM64_INSTR_PT(545) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011011"));
MQQ546:ROM64_INSTR_PT(546) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011011"));
MQQ547:ROM64_INSTR_PT(547) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ548:ROM64_INSTR_PT(548) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111011"));
MQQ549:ROM64_INSTR_PT(549) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101011"));
MQQ550:ROM64_INSTR_PT(550) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011011"));
MQQ551:ROM64_INSTR_PT(551) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ552:ROM64_INSTR_PT(552) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100011"));
MQQ553:ROM64_INSTR_PT(553) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100011"));
MQQ554:ROM64_INSTR_PT(554) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010011"));
MQQ555:ROM64_INSTR_PT(555) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110011"));
MQQ556:ROM64_INSTR_PT(556) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001011"));
MQQ557:ROM64_INSTR_PT(557) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101011"));
MQQ558:ROM64_INSTR_PT(558) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011011"));
MQQ559:ROM64_INSTR_PT(559) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011011"));
MQQ560:ROM64_INSTR_PT(560) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111011"));
MQQ561:ROM64_INSTR_PT(561) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101011"));
MQQ562:ROM64_INSTR_PT(562) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011011"));
MQQ563:ROM64_INSTR_PT(563) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111011"));
MQQ564:ROM64_INSTR_PT(564) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111011"));
MQQ565:ROM64_INSTR_PT(565) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ566:ROM64_INSTR_PT(566) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000111"));
MQQ567:ROM64_INSTR_PT(567) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000111"));
MQQ568:ROM64_INSTR_PT(568) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110000111"));
MQQ569:ROM64_INSTR_PT(569) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000111"));
MQQ570:ROM64_INSTR_PT(570) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000111"));
MQQ571:ROM64_INSTR_PT(571) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000111"));
MQQ572:ROM64_INSTR_PT(572) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010100111"));
MQQ573:ROM64_INSTR_PT(573) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100111"));
MQQ574:ROM64_INSTR_PT(574) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100111"));
MQQ575:ROM64_INSTR_PT(575) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100111"));
MQQ576:ROM64_INSTR_PT(576) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100111"));
MQQ577:ROM64_INSTR_PT(577) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100111"));
MQQ578:ROM64_INSTR_PT(578) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000111"));
MQQ579:ROM64_INSTR_PT(579) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010111"));
MQQ580:ROM64_INSTR_PT(580) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010111"));
MQQ581:ROM64_INSTR_PT(581) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001010111"));
MQQ582:ROM64_INSTR_PT(582) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010111"));
MQQ583:ROM64_INSTR_PT(583) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110111"));
MQQ584:ROM64_INSTR_PT(584) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010111"));
MQQ585:ROM64_INSTR_PT(585) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000111"));
MQQ586:ROM64_INSTR_PT(586) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100111"));
MQQ587:ROM64_INSTR_PT(587) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010111"));
MQQ588:ROM64_INSTR_PT(588) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001111"));
MQQ589:ROM64_INSTR_PT(589) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100001111"));
MQQ590:ROM64_INSTR_PT(590) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001111"));
MQQ591:ROM64_INSTR_PT(591) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001111"));
MQQ592:ROM64_INSTR_PT(592) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001111"));
MQQ593:ROM64_INSTR_PT(593) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001111"));
MQQ594:ROM64_INSTR_PT(594) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001111"));
MQQ595:ROM64_INSTR_PT(595) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000101111"));
MQQ596:ROM64_INSTR_PT(596) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010101111"));
MQQ597:ROM64_INSTR_PT(597) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001101111"));
MQQ598:ROM64_INSTR_PT(598) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101111"));
MQQ599:ROM64_INSTR_PT(599) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101111"));
MQQ600:ROM64_INSTR_PT(600) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101111"));
MQQ601:ROM64_INSTR_PT(601) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011111"));
MQQ602:ROM64_INSTR_PT(602) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011111"));
MQQ603:ROM64_INSTR_PT(603) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001011111"));
MQQ604:ROM64_INSTR_PT(604) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111111"));
MQQ605:ROM64_INSTR_PT(605) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111111"));
MQQ606:ROM64_INSTR_PT(606) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111111"));
MQQ607:ROM64_INSTR_PT(607) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ608:ROM64_INSTR_PT(608) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011111"));
MQQ609:ROM64_INSTR_PT(609) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ610:ROM64_INSTR_PT(610) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111111"));
MQQ611:ROM64_INSTR_PT(611) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111111"));
MQQ612:ROM64_INSTR_PT(612) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111111"));
MQQ613:ROM64_INSTR_PT(613) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101111"));
MQQ614:ROM64_INSTR_PT(614) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ615:ROM64_INSTR_PT(615) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111111"));
MQQ616:ROM64_INSTR_PT(616) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111111"));
MQQ617:ROM64_INSTR_PT(617) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ618:ROM64_INSTR_PT(618) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ619:ROM64_INSTR_PT(619) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110111"));
MQQ620:ROM64_INSTR_PT(620) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100111"));
MQQ621:ROM64_INSTR_PT(621) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011111"));
MQQ622:ROM64_INSTR_PT(622) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ623:ROM64_INSTR_PT(623) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111111"));
MQQ624:ROM64_INSTR_PT(624) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ625:ROM64_INSTR_PT(625) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ626:ROM64_INSTR_PT(626) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001111"));
MQQ627:ROM64_INSTR_PT(627) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ628:ROM64_INSTR_PT(628) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ629:ROM64_INSTR_PT(629) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ630:ROM64_INSTR_PT(630) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ631:ROM64_INSTR_PT(631) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110011"));
MQQ632:ROM64_INSTR_PT(632) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101011"));
MQQ633:ROM64_INSTR_PT(633) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011011"));
MQQ634:ROM64_INSTR_PT(634) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111011"));
MQQ635:ROM64_INSTR_PT(635) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111011"));
MQQ636:ROM64_INSTR_PT(636) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ637:ROM64_INSTR_PT(637) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ638:ROM64_INSTR_PT(638) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("10011"));
MQQ639:ROM64_INSTR_PT(639) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100111"));
MQQ640:ROM64_INSTR_PT(640) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110111"));
MQQ641:ROM64_INSTR_PT(641) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000111"));
MQQ642:ROM64_INSTR_PT(642) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ643:ROM64_INSTR_PT(643) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ644:ROM64_INSTR_PT(644) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ645:ROM64_INSTR_PT(645) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110111"));
MQQ646:ROM64_INSTR_PT(646) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011111"));
MQQ647:ROM64_INSTR_PT(647) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ648:ROM64_INSTR_PT(648) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ649:ROM64_INSTR_PT(649) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ650:ROM64_INSTR_PT(650) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ651:ROM64_INSTR_PT(651) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("10111"));
MQQ652:ROM64_INSTR_PT(652) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ653:ROM64_INSTR_PT(653) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ654:ROM64_INSTR_PT(654) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000001"));
MQQ655:ROM64_INSTR_PT(655) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110001"));
MQQ656:ROM64_INSTR_PT(656) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110001"));
MQQ657:ROM64_INSTR_PT(657) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101001"));
MQQ658:ROM64_INSTR_PT(658) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001001"));
MQQ659:ROM64_INSTR_PT(659) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011001"));
MQQ660:ROM64_INSTR_PT(660) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101001"));
MQQ661:ROM64_INSTR_PT(661) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000101"));
MQQ662:ROM64_INSTR_PT(662) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000101"));
MQQ663:ROM64_INSTR_PT(663) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100101"));
MQQ664:ROM64_INSTR_PT(664) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110101"));
MQQ665:ROM64_INSTR_PT(665) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001101"));
MQQ666:ROM64_INSTR_PT(666) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011101"));
MQQ667:ROM64_INSTR_PT(667) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011101"));
MQQ668:ROM64_INSTR_PT(668) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000001"));
MQQ669:ROM64_INSTR_PT(669) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010001"));
MQQ670:ROM64_INSTR_PT(670) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110001"));
MQQ671:ROM64_INSTR_PT(671) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001001"));
MQQ672:ROM64_INSTR_PT(672) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0010101"));
MQQ673:ROM64_INSTR_PT(673) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011101"));
MQQ674:ROM64_INSTR_PT(674) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000011"));
MQQ675:ROM64_INSTR_PT(675) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100011"));
MQQ676:ROM64_INSTR_PT(676) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ677:ROM64_INSTR_PT(677) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ678:ROM64_INSTR_PT(678) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101011"));
MQQ679:ROM64_INSTR_PT(679) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011011"));
MQQ680:ROM64_INSTR_PT(680) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011011"));
MQQ681:ROM64_INSTR_PT(681) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ682:ROM64_INSTR_PT(682) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ683:ROM64_INSTR_PT(683) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010011"));
MQQ684:ROM64_INSTR_PT(684) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100111"));
MQQ685:ROM64_INSTR_PT(685) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010111"));
MQQ686:ROM64_INSTR_PT(686) <=
    Eq(( ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0111"));
MQQ687:ROM64_INSTR_PT(687) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001111"));
MQQ688:ROM64_INSTR_PT(688) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101111"));
MQQ689:ROM64_INSTR_PT(689) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011111"));
MQQ690:ROM64_INSTR_PT(690) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ691:ROM64_INSTR_PT(691) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ692:ROM64_INSTR_PT(692) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101111"));
MQQ693:ROM64_INSTR_PT(693) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ694:ROM64_INSTR_PT(694) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000111"));
MQQ695:ROM64_INSTR_PT(695) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110111"));
MQQ696:ROM64_INSTR_PT(696) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("000111"));
MQQ697:ROM64_INSTR_PT(697) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ698:ROM64_INSTR_PT(698) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011111"));
MQQ699:ROM64_INSTR_PT(699) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ700:ROM64_INSTR_PT(700) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011011"));
MQQ701:ROM64_INSTR_PT(701) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ702:ROM64_INSTR_PT(702) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ703:ROM64_INSTR_PT(703) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101111"));
MQQ704:ROM64_INSTR_PT(704) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ705:ROM64_INSTR_PT(705) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ706:ROM64_INSTR_PT(706) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000001"));
MQQ707:ROM64_INSTR_PT(707) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010001"));
MQQ708:ROM64_INSTR_PT(708) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001001"));
MQQ709:ROM64_INSTR_PT(709) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111001"));
MQQ710:ROM64_INSTR_PT(710) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100101"));
MQQ711:ROM64_INSTR_PT(711) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100001"));
MQQ712:ROM64_INSTR_PT(712) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111101"));
MQQ713:ROM64_INSTR_PT(713) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0110111"));
MQQ714:ROM64_INSTR_PT(714) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ715:ROM64_INSTR_PT(715) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ716:ROM64_INSTR_PT(716) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ717:ROM64_INSTR_PT(717) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011111"));
MQQ718:ROM64_INSTR_PT(718) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ719:ROM64_INSTR_PT(719) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100101"));
MQQ720:ROM64_INSTR_PT(720) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ721:ROM64_INSTR_PT(721) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101"));
MQQ722:ROM64_INSTR_PT(722) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100000"));
MQQ723:ROM64_INSTR_PT(723) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100000"));
MQQ724:ROM64_INSTR_PT(724) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("010010000"));
MQQ725:ROM64_INSTR_PT(725) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000110000"));
MQQ726:ROM64_INSTR_PT(726) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ727:ROM64_INSTR_PT(727) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100000"));
MQQ728:ROM64_INSTR_PT(728) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("010001000"));
MQQ729:ROM64_INSTR_PT(729) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11011000"));
MQQ730:ROM64_INSTR_PT(730) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111000"));
MQQ731:ROM64_INSTR_PT(731) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0111000"));
MQQ732:ROM64_INSTR_PT(732) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110000"));
MQQ733:ROM64_INSTR_PT(733) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00000100"));
MQQ734:ROM64_INSTR_PT(734) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000100"));
MQQ735:ROM64_INSTR_PT(735) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100100"));
MQQ736:ROM64_INSTR_PT(736) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1100100"));
MQQ737:ROM64_INSTR_PT(737) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100100"));
MQQ738:ROM64_INSTR_PT(738) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("010010100"));
MQQ739:ROM64_INSTR_PT(739) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ740:ROM64_INSTR_PT(740) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ741:ROM64_INSTR_PT(741) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("10011100"));
MQQ742:ROM64_INSTR_PT(742) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101100"));
MQQ743:ROM64_INSTR_PT(743) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0111100"));
MQQ744:ROM64_INSTR_PT(744) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100100"));
MQQ745:ROM64_INSTR_PT(745) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100000"));
MQQ746:ROM64_INSTR_PT(746) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1100000"));
MQQ747:ROM64_INSTR_PT(747) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00000100"));
MQQ748:ROM64_INSTR_PT(748) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0101100"));
MQQ749:ROM64_INSTR_PT(749) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011100"));
MQQ750:ROM64_INSTR_PT(750) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ751:ROM64_INSTR_PT(751) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11100"));
MQQ752:ROM64_INSTR_PT(752) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000"));
MQQ753:ROM64_INSTR_PT(753) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100010"));
MQQ754:ROM64_INSTR_PT(754) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00010010"));
MQQ755:ROM64_INSTR_PT(755) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00000010"));
MQQ756:ROM64_INSTR_PT(756) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11001010"));
MQQ757:ROM64_INSTR_PT(757) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111010"));
MQQ758:ROM64_INSTR_PT(758) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1111010"));
MQQ759:ROM64_INSTR_PT(759) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101010"));
MQQ760:ROM64_INSTR_PT(760) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1000110"));
MQQ761:ROM64_INSTR_PT(761) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("110100110"));
MQQ762:ROM64_INSTR_PT(762) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0010110"));
MQQ763:ROM64_INSTR_PT(763) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("010110"));
MQQ764:ROM64_INSTR_PT(764) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0001110"));
MQQ765:ROM64_INSTR_PT(765) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011110"));
MQQ766:ROM64_INSTR_PT(766) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("10011110"));
MQQ767:ROM64_INSTR_PT(767) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ768:ROM64_INSTR_PT(768) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("0110"));
MQQ769:ROM64_INSTR_PT(769) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011110"));
MQQ770:ROM64_INSTR_PT(770) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ771:ROM64_INSTR_PT(771) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("010110"));
MQQ772:ROM64_INSTR_PT(772) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("10000"));
MQQ773:ROM64_INSTR_PT(773) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ774:ROM64_INSTR_PT(774) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011100"));
MQQ775:ROM64_INSTR_PT(775) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("00100"));
MQQ776:ROM64_INSTR_PT(776) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100010"));
MQQ777:ROM64_INSTR_PT(777) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11010010"));
MQQ778:ROM64_INSTR_PT(778) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101010"));
MQQ779:ROM64_INSTR_PT(779) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01110"));
MQQ780:ROM64_INSTR_PT(780) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01110"));
MQQ781:ROM64_INSTR_PT(781) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01000001"));
MQQ782:ROM64_INSTR_PT(782) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("110100001"));
MQQ783:ROM64_INSTR_PT(783) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01010001"));
MQQ784:ROM64_INSTR_PT(784) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11010001"));
MQQ785:ROM64_INSTR_PT(785) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1010001"));
MQQ786:ROM64_INSTR_PT(786) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000001"));
MQQ787:ROM64_INSTR_PT(787) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("010001"));
MQQ788:ROM64_INSTR_PT(788) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0001001"));
MQQ789:ROM64_INSTR_PT(789) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("001001"));
MQQ790:ROM64_INSTR_PT(790) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011001"));
MQQ791:ROM64_INSTR_PT(791) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111001"));
MQQ792:ROM64_INSTR_PT(792) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011001"));
MQQ793:ROM64_INSTR_PT(793) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111001"));
MQQ794:ROM64_INSTR_PT(794) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00100101"));
MQQ795:ROM64_INSTR_PT(795) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00010101"));
MQQ796:ROM64_INSTR_PT(796) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011101"));
MQQ797:ROM64_INSTR_PT(797) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("10011101"));
MQQ798:ROM64_INSTR_PT(798) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110101"));
MQQ799:ROM64_INSTR_PT(799) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("10101"));
MQQ800:ROM64_INSTR_PT(800) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11101"));
MQQ801:ROM64_INSTR_PT(801) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000101"));
MQQ802:ROM64_INSTR_PT(802) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000101"));
MQQ803:ROM64_INSTR_PT(803) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11101"));
MQQ804:ROM64_INSTR_PT(804) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000100011"));
MQQ805:ROM64_INSTR_PT(805) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01110011"));
MQQ806:ROM64_INSTR_PT(806) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00000011"));
MQQ807:ROM64_INSTR_PT(807) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000011"));
MQQ808:ROM64_INSTR_PT(808) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000011"));
MQQ809:ROM64_INSTR_PT(809) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1010011"));
MQQ810:ROM64_INSTR_PT(810) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("010011"));
MQQ811:ROM64_INSTR_PT(811) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01101011"));
MQQ812:ROM64_INSTR_PT(812) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00001011"));
MQQ813:ROM64_INSTR_PT(813) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ814:ROM64_INSTR_PT(814) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101011"));
MQQ815:ROM64_INSTR_PT(815) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ816:ROM64_INSTR_PT(816) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100111"));
MQQ817:ROM64_INSTR_PT(817) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00010111"));
MQQ818:ROM64_INSTR_PT(818) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ819:ROM64_INSTR_PT(819) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1110111"));
MQQ820:ROM64_INSTR_PT(820) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11010111"));
MQQ821:ROM64_INSTR_PT(821) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000101111"));
MQQ822:ROM64_INSTR_PT(822) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01101111"));
MQQ823:ROM64_INSTR_PT(823) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ824:ROM64_INSTR_PT(824) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ825:ROM64_INSTR_PT(825) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ826:ROM64_INSTR_PT(826) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ827:ROM64_INSTR_PT(827) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101011"));
MQQ828:ROM64_INSTR_PT(828) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0110111"));
MQQ829:ROM64_INSTR_PT(829) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ830:ROM64_INSTR_PT(830) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ831:ROM64_INSTR_PT(831) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("0111"));
MQQ832:ROM64_INSTR_PT(832) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ833:ROM64_INSTR_PT(833) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ834:ROM64_INSTR_PT(834) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110001"));
MQQ835:ROM64_INSTR_PT(835) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1001101"));
MQQ836:ROM64_INSTR_PT(836) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101101"));
MQQ837:ROM64_INSTR_PT(837) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101011"));
MQQ838:ROM64_INSTR_PT(838) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1111011"));
MQQ839:ROM64_INSTR_PT(839) <=
    Eq(( ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("011"));
MQQ840:ROM64_INSTR_PT(840) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000111"));
MQQ841:ROM64_INSTR_PT(841) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ842:ROM64_INSTR_PT(842) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101111"));
MQQ843:ROM64_INSTR_PT(843) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01111"));
MQQ844:ROM64_INSTR_PT(844) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ845:ROM64_INSTR_PT(845) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ846:ROM64_INSTR_PT(846) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011111"));
MQQ847:ROM64_INSTR_PT(847) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("000101"));
MQQ848:ROM64_INSTR_PT(848) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01101"));
MQQ849:ROM64_INSTR_PT(849) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ850:ROM64_INSTR_PT(850) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("1111"));
MQQ851:ROM64_INSTR_PT(851) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01001"));
MQQ852:ROM64_INSTR_PT(852) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1001000"));
MQQ853:ROM64_INSTR_PT(853) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("110000"));
MQQ854:ROM64_INSTR_PT(854) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("00011100"));
MQQ855:ROM64_INSTR_PT(855) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("00000010"));
MQQ856:ROM64_INSTR_PT(856) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0100010"));
MQQ857:ROM64_INSTR_PT(857) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0000010"));
MQQ858:ROM64_INSTR_PT(858) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("101110"));
MQQ859:ROM64_INSTR_PT(859) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1101110"));
MQQ860:ROM64_INSTR_PT(860) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("000110"));
MQQ861:ROM64_INSTR_PT(861) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1001100"));
MQQ862:ROM64_INSTR_PT(862) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("1110"));
MQQ863:ROM64_INSTR_PT(863) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("010"));
MQQ864:ROM64_INSTR_PT(864) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0100101"));
MQQ865:ROM64_INSTR_PT(865) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1100101"));
MQQ866:ROM64_INSTR_PT(866) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1001101"));
MQQ867:ROM64_INSTR_PT(867) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1101101"));
MQQ868:ROM64_INSTR_PT(868) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("01011"));
MQQ869:ROM64_INSTR_PT(869) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ870:ROM64_INSTR_PT(870) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0011111"));
MQQ871:ROM64_INSTR_PT(871) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("100111"));
MQQ872:ROM64_INSTR_PT(872) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ873:ROM64_INSTR_PT(873) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ874:ROM64_INSTR_PT(874) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ875:ROM64_INSTR_PT(875) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("01111"));
MQQ876:ROM64_INSTR_PT(876) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("101"));
MQQ877:ROM64_INSTR_PT(877) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("010001"));
MQQ878:ROM64_INSTR_PT(878) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("01111"));
MQQ879:ROM64_INSTR_PT(879) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("111"));
MQQ880:ROM64_INSTR_PT(880) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) ) , STD_ULOGIC_VECTOR'("01110"));
MQQ881:ROM64_INSTR_PT(881) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(6)
     ) , STD_ULOGIC_VECTOR'("00"));
MQQ882:ROM64_INSTR_PT(882) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) ) , STD_ULOGIC_VECTOR'("111"));
MQQ883:ROM64_INSTR_PT(883) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ884:ROM64_INSTR_PT(884) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5)
     ) , STD_ULOGIC_VECTOR'("00"));
MQQ885:ROM64_INSTR_PT(885) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) ) , STD_ULOGIC_VECTOR'("111"));
MQQ886:ROM64_INSTR_PT(886) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) ) , STD_ULOGIC_VECTOR'("111"));
MQQ887:ROM64_INSTR_PT(887) <=
    Eq(( ROM_ADDR_L2(2) ) , STD_ULOGIC'('1'));
MQQ888:ROM64_INSTR_PT(888) <=
    Eq(( ROM_ADDR_L2(1) ) , STD_ULOGIC'('1'));
MQQ889:ROM64_INSTR_PT(889) <=
    Eq(( ROM_ADDR_L2(0) ) , STD_ULOGIC'('0'));
MQQ890:ROM64_INSTR_PT(890) <=
    '1';
-- Table ROM64_INSTR Signal Assignments for Outputs
MQQ891:TEMPLATE(0) <= 
    (ROM64_INSTR_PT(29) OR ROM64_INSTR_PT(35)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(65)
     OR ROM64_INSTR_PT(74) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(112) OR ROM64_INSTR_PT(119)
     OR ROM64_INSTR_PT(129) OR ROM64_INSTR_PT(134)
     OR ROM64_INSTR_PT(143) OR ROM64_INSTR_PT(158)
     OR ROM64_INSTR_PT(160) OR ROM64_INSTR_PT(176)
     OR ROM64_INSTR_PT(177) OR ROM64_INSTR_PT(179)
     OR ROM64_INSTR_PT(183) OR ROM64_INSTR_PT(221)
     OR ROM64_INSTR_PT(225) OR ROM64_INSTR_PT(233)
     OR ROM64_INSTR_PT(237) OR ROM64_INSTR_PT(242)
     OR ROM64_INSTR_PT(259) OR ROM64_INSTR_PT(294)
     OR ROM64_INSTR_PT(296) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(339) OR ROM64_INSTR_PT(350)
     OR ROM64_INSTR_PT(354) OR ROM64_INSTR_PT(355)
     OR ROM64_INSTR_PT(358) OR ROM64_INSTR_PT(359)
     OR ROM64_INSTR_PT(362) OR ROM64_INSTR_PT(367)
     OR ROM64_INSTR_PT(368) OR ROM64_INSTR_PT(378)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(389)
     OR ROM64_INSTR_PT(392) OR ROM64_INSTR_PT(402)
     OR ROM64_INSTR_PT(428) OR ROM64_INSTR_PT(435)
     OR ROM64_INSTR_PT(470) OR ROM64_INSTR_PT(477)
     OR ROM64_INSTR_PT(527) OR ROM64_INSTR_PT(557)
     OR ROM64_INSTR_PT(564) OR ROM64_INSTR_PT(572)
     OR ROM64_INSTR_PT(590) OR ROM64_INSTR_PT(602)
     OR ROM64_INSTR_PT(610) OR ROM64_INSTR_PT(619)
     OR ROM64_INSTR_PT(653) OR ROM64_INSTR_PT(657)
     OR ROM64_INSTR_PT(664) OR ROM64_INSTR_PT(694)
     OR ROM64_INSTR_PT(695) OR ROM64_INSTR_PT(702)
     OR ROM64_INSTR_PT(716) OR ROM64_INSTR_PT(719)
     OR ROM64_INSTR_PT(720) OR ROM64_INSTR_PT(721)
     OR ROM64_INSTR_PT(736) OR ROM64_INSTR_PT(770)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(832)
     OR ROM64_INSTR_PT(834) OR ROM64_INSTR_PT(858)
     OR ROM64_INSTR_PT(873));
MQQ892:TEMPLATE(1) <= 
    (ROM64_INSTR_PT(2) OR ROM64_INSTR_PT(4)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(8)
     OR ROM64_INSTR_PT(9) OR ROM64_INSTR_PT(10)
     OR ROM64_INSTR_PT(11) OR ROM64_INSTR_PT(14)
     OR ROM64_INSTR_PT(15) OR ROM64_INSTR_PT(17)
     OR ROM64_INSTR_PT(18) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(25)
     OR ROM64_INSTR_PT(34) OR ROM64_INSTR_PT(36)
     OR ROM64_INSTR_PT(38) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(43)
     OR ROM64_INSTR_PT(49) OR ROM64_INSTR_PT(51)
     OR ROM64_INSTR_PT(52) OR ROM64_INSTR_PT(53)
     OR ROM64_INSTR_PT(55) OR ROM64_INSTR_PT(56)
     OR ROM64_INSTR_PT(61) OR ROM64_INSTR_PT(64)
     OR ROM64_INSTR_PT(68) OR ROM64_INSTR_PT(69)
     OR ROM64_INSTR_PT(70) OR ROM64_INSTR_PT(71)
     OR ROM64_INSTR_PT(73) OR ROM64_INSTR_PT(75)
     OR ROM64_INSTR_PT(77) OR ROM64_INSTR_PT(78)
     OR ROM64_INSTR_PT(82) OR ROM64_INSTR_PT(83)
     OR ROM64_INSTR_PT(86) OR ROM64_INSTR_PT(89)
     OR ROM64_INSTR_PT(90) OR ROM64_INSTR_PT(92)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(95)
     OR ROM64_INSTR_PT(96) OR ROM64_INSTR_PT(97)
     OR ROM64_INSTR_PT(99) OR ROM64_INSTR_PT(100)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(102)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(105)
     OR ROM64_INSTR_PT(106) OR ROM64_INSTR_PT(108)
     OR ROM64_INSTR_PT(109) OR ROM64_INSTR_PT(110)
     OR ROM64_INSTR_PT(113) OR ROM64_INSTR_PT(116)
     OR ROM64_INSTR_PT(117) OR ROM64_INSTR_PT(118)
     OR ROM64_INSTR_PT(124) OR ROM64_INSTR_PT(127)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(144)
     OR ROM64_INSTR_PT(145) OR ROM64_INSTR_PT(148)
     OR ROM64_INSTR_PT(153) OR ROM64_INSTR_PT(161)
     OR ROM64_INSTR_PT(162) OR ROM64_INSTR_PT(164)
     OR ROM64_INSTR_PT(169) OR ROM64_INSTR_PT(170)
     OR ROM64_INSTR_PT(171) OR ROM64_INSTR_PT(172)
     OR ROM64_INSTR_PT(173) OR ROM64_INSTR_PT(175)
     OR ROM64_INSTR_PT(180) OR ROM64_INSTR_PT(184)
     OR ROM64_INSTR_PT(185) OR ROM64_INSTR_PT(186)
     OR ROM64_INSTR_PT(188) OR ROM64_INSTR_PT(193)
     OR ROM64_INSTR_PT(195) OR ROM64_INSTR_PT(196)
     OR ROM64_INSTR_PT(199) OR ROM64_INSTR_PT(201)
     OR ROM64_INSTR_PT(202) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(205) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(208) OR ROM64_INSTR_PT(214)
     OR ROM64_INSTR_PT(215) OR ROM64_INSTR_PT(216)
     OR ROM64_INSTR_PT(217) OR ROM64_INSTR_PT(218)
     OR ROM64_INSTR_PT(222) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(226) OR ROM64_INSTR_PT(229)
     OR ROM64_INSTR_PT(230) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(241) OR ROM64_INSTR_PT(243)
     OR ROM64_INSTR_PT(244) OR ROM64_INSTR_PT(252)
     OR ROM64_INSTR_PT(254) OR ROM64_INSTR_PT(257)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(263)
     OR ROM64_INSTR_PT(264) OR ROM64_INSTR_PT(265)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(269)
     OR ROM64_INSTR_PT(270) OR ROM64_INSTR_PT(271)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(275)
     OR ROM64_INSTR_PT(276) OR ROM64_INSTR_PT(277)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(282)
     OR ROM64_INSTR_PT(284) OR ROM64_INSTR_PT(285)
     OR ROM64_INSTR_PT(286) OR ROM64_INSTR_PT(287)
     OR ROM64_INSTR_PT(292) OR ROM64_INSTR_PT(293)
     OR ROM64_INSTR_PT(297) OR ROM64_INSTR_PT(298)
     OR ROM64_INSTR_PT(299) OR ROM64_INSTR_PT(302)
     OR ROM64_INSTR_PT(305) OR ROM64_INSTR_PT(308)
     OR ROM64_INSTR_PT(315) OR ROM64_INSTR_PT(322)
     OR ROM64_INSTR_PT(325) OR ROM64_INSTR_PT(331)
     OR ROM64_INSTR_PT(333) OR ROM64_INSTR_PT(345)
     OR ROM64_INSTR_PT(349) OR ROM64_INSTR_PT(351)
     OR ROM64_INSTR_PT(357) OR ROM64_INSTR_PT(364)
     OR ROM64_INSTR_PT(365) OR ROM64_INSTR_PT(366)
     OR ROM64_INSTR_PT(369) OR ROM64_INSTR_PT(371)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(375)
     OR ROM64_INSTR_PT(377) OR ROM64_INSTR_PT(379)
     OR ROM64_INSTR_PT(381) OR ROM64_INSTR_PT(383)
     OR ROM64_INSTR_PT(385) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(391) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(403) OR ROM64_INSTR_PT(404)
     OR ROM64_INSTR_PT(405) OR ROM64_INSTR_PT(408)
     OR ROM64_INSTR_PT(409) OR ROM64_INSTR_PT(410)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(419) OR ROM64_INSTR_PT(420)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(424)
     OR ROM64_INSTR_PT(425) OR ROM64_INSTR_PT(426)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(429)
     OR ROM64_INSTR_PT(430) OR ROM64_INSTR_PT(432)
     OR ROM64_INSTR_PT(433) OR ROM64_INSTR_PT(434)
     OR ROM64_INSTR_PT(437) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(439) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(443) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(451)
     OR ROM64_INSTR_PT(453) OR ROM64_INSTR_PT(454)
     OR ROM64_INSTR_PT(455) OR ROM64_INSTR_PT(456)
     OR ROM64_INSTR_PT(457) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(460) OR ROM64_INSTR_PT(463)
     OR ROM64_INSTR_PT(466) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(478) OR ROM64_INSTR_PT(480)
     OR ROM64_INSTR_PT(481) OR ROM64_INSTR_PT(482)
     OR ROM64_INSTR_PT(483) OR ROM64_INSTR_PT(484)
     OR ROM64_INSTR_PT(485) OR ROM64_INSTR_PT(490)
     OR ROM64_INSTR_PT(493) OR ROM64_INSTR_PT(495)
     OR ROM64_INSTR_PT(497) OR ROM64_INSTR_PT(498)
     OR ROM64_INSTR_PT(499) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(505)
     OR ROM64_INSTR_PT(506) OR ROM64_INSTR_PT(508)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(510)
     OR ROM64_INSTR_PT(511) OR ROM64_INSTR_PT(512)
     OR ROM64_INSTR_PT(514) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(521) OR ROM64_INSTR_PT(522)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(525)
     OR ROM64_INSTR_PT(530) OR ROM64_INSTR_PT(531)
     OR ROM64_INSTR_PT(532) OR ROM64_INSTR_PT(534)
     OR ROM64_INSTR_PT(535) OR ROM64_INSTR_PT(536)
     OR ROM64_INSTR_PT(537) OR ROM64_INSTR_PT(539)
     OR ROM64_INSTR_PT(540) OR ROM64_INSTR_PT(542)
     OR ROM64_INSTR_PT(544) OR ROM64_INSTR_PT(545)
     OR ROM64_INSTR_PT(546) OR ROM64_INSTR_PT(548)
     OR ROM64_INSTR_PT(549) OR ROM64_INSTR_PT(552)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(555) OR ROM64_INSTR_PT(558)
     OR ROM64_INSTR_PT(559) OR ROM64_INSTR_PT(563)
     OR ROM64_INSTR_PT(566) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(569) OR ROM64_INSTR_PT(570)
     OR ROM64_INSTR_PT(571) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(577)
     OR ROM64_INSTR_PT(579) OR ROM64_INSTR_PT(580)
     OR ROM64_INSTR_PT(581) OR ROM64_INSTR_PT(582)
     OR ROM64_INSTR_PT(583) OR ROM64_INSTR_PT(584)
     OR ROM64_INSTR_PT(586) OR ROM64_INSTR_PT(588)
     OR ROM64_INSTR_PT(589) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(592) OR ROM64_INSTR_PT(593)
     OR ROM64_INSTR_PT(595) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(598) OR ROM64_INSTR_PT(599)
     OR ROM64_INSTR_PT(600) OR ROM64_INSTR_PT(603)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(606)
     OR ROM64_INSTR_PT(607) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(611) OR ROM64_INSTR_PT(612)
     OR ROM64_INSTR_PT(613) OR ROM64_INSTR_PT(614)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(616)
     OR ROM64_INSTR_PT(617) OR ROM64_INSTR_PT(618)
     OR ROM64_INSTR_PT(623) OR ROM64_INSTR_PT(626)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(629) OR ROM64_INSTR_PT(633)
     OR ROM64_INSTR_PT(637) OR ROM64_INSTR_PT(639)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(643)
     OR ROM64_INSTR_PT(644) OR ROM64_INSTR_PT(646)
     OR ROM64_INSTR_PT(655) OR ROM64_INSTR_PT(660)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(666)
     OR ROM64_INSTR_PT(678) OR ROM64_INSTR_PT(679)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(682)
     OR ROM64_INSTR_PT(687) OR ROM64_INSTR_PT(703)
     OR ROM64_INSTR_PT(713) OR ROM64_INSTR_PT(717)
     OR ROM64_INSTR_PT(722) OR ROM64_INSTR_PT(731)
     OR ROM64_INSTR_PT(741) OR ROM64_INSTR_PT(744)
     OR ROM64_INSTR_PT(753) OR ROM64_INSTR_PT(761)
     OR ROM64_INSTR_PT(769) OR ROM64_INSTR_PT(776)
     OR ROM64_INSTR_PT(791) OR ROM64_INSTR_PT(801)
     OR ROM64_INSTR_PT(808) OR ROM64_INSTR_PT(811)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(822)
     OR ROM64_INSTR_PT(824) OR ROM64_INSTR_PT(846)
     OR ROM64_INSTR_PT(849) OR ROM64_INSTR_PT(852)
     OR ROM64_INSTR_PT(854) OR ROM64_INSTR_PT(855)
     OR ROM64_INSTR_PT(856) OR ROM64_INSTR_PT(864)
     OR ROM64_INSTR_PT(869) OR ROM64_INSTR_PT(870)
     OR ROM64_INSTR_PT(872) OR ROM64_INSTR_PT(886)
    );
MQQ893:TEMPLATE(2) <= 
    (ROM64_INSTR_PT(2) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(10)
     OR ROM64_INSTR_PT(14) OR ROM64_INSTR_PT(15)
     OR ROM64_INSTR_PT(18) OR ROM64_INSTR_PT(20)
     OR ROM64_INSTR_PT(25) OR ROM64_INSTR_PT(28)
     OR ROM64_INSTR_PT(33) OR ROM64_INSTR_PT(36)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(43)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(56)
     OR ROM64_INSTR_PT(60) OR ROM64_INSTR_PT(66)
     OR ROM64_INSTR_PT(69) OR ROM64_INSTR_PT(73)
     OR ROM64_INSTR_PT(77) OR ROM64_INSTR_PT(78)
     OR ROM64_INSTR_PT(79) OR ROM64_INSTR_PT(82)
     OR ROM64_INSTR_PT(89) OR ROM64_INSTR_PT(92)
     OR ROM64_INSTR_PT(95) OR ROM64_INSTR_PT(96)
     OR ROM64_INSTR_PT(97) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(104)
     OR ROM64_INSTR_PT(106) OR ROM64_INSTR_PT(108)
     OR ROM64_INSTR_PT(109) OR ROM64_INSTR_PT(110)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(124)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(142)
     OR ROM64_INSTR_PT(145) OR ROM64_INSTR_PT(146)
     OR ROM64_INSTR_PT(147) OR ROM64_INSTR_PT(150)
     OR ROM64_INSTR_PT(151) OR ROM64_INSTR_PT(153)
     OR ROM64_INSTR_PT(161) OR ROM64_INSTR_PT(166)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(172)
     OR ROM64_INSTR_PT(173) OR ROM64_INSTR_PT(174)
     OR ROM64_INSTR_PT(175) OR ROM64_INSTR_PT(184)
     OR ROM64_INSTR_PT(187) OR ROM64_INSTR_PT(188)
     OR ROM64_INSTR_PT(190) OR ROM64_INSTR_PT(191)
     OR ROM64_INSTR_PT(193) OR ROM64_INSTR_PT(195)
     OR ROM64_INSTR_PT(202) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(205) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(207) OR ROM64_INSTR_PT(208)
     OR ROM64_INSTR_PT(209) OR ROM64_INSTR_PT(216)
     OR ROM64_INSTR_PT(219) OR ROM64_INSTR_PT(228)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(231) OR ROM64_INSTR_PT(240)
     OR ROM64_INSTR_PT(243) OR ROM64_INSTR_PT(247)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(254)
     OR ROM64_INSTR_PT(257) OR ROM64_INSTR_PT(258)
     OR ROM64_INSTR_PT(260) OR ROM64_INSTR_PT(261)
     OR ROM64_INSTR_PT(265) OR ROM64_INSTR_PT(269)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(277)
     OR ROM64_INSTR_PT(281) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(288) OR ROM64_INSTR_PT(292)
     OR ROM64_INSTR_PT(295) OR ROM64_INSTR_PT(304)
     OR ROM64_INSTR_PT(307) OR ROM64_INSTR_PT(309)
     OR ROM64_INSTR_PT(313) OR ROM64_INSTR_PT(324)
     OR ROM64_INSTR_PT(325) OR ROM64_INSTR_PT(327)
     OR ROM64_INSTR_PT(332) OR ROM64_INSTR_PT(333)
     OR ROM64_INSTR_PT(334) OR ROM64_INSTR_PT(340)
     OR ROM64_INSTR_PT(341) OR ROM64_INSTR_PT(342)
     OR ROM64_INSTR_PT(345) OR ROM64_INSTR_PT(351)
     OR ROM64_INSTR_PT(352) OR ROM64_INSTR_PT(357)
     OR ROM64_INSTR_PT(361) OR ROM64_INSTR_PT(365)
     OR ROM64_INSTR_PT(366) OR ROM64_INSTR_PT(369)
     OR ROM64_INSTR_PT(371) OR ROM64_INSTR_PT(372)
     OR ROM64_INSTR_PT(374) OR ROM64_INSTR_PT(377)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(388) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(396)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(403)
     OR ROM64_INSTR_PT(405) OR ROM64_INSTR_PT(406)
     OR ROM64_INSTR_PT(408) OR ROM64_INSTR_PT(409)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(419) OR ROM64_INSTR_PT(420)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(425)
     OR ROM64_INSTR_PT(426) OR ROM64_INSTR_PT(429)
     OR ROM64_INSTR_PT(430) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(439) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(443) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(448)
     OR ROM64_INSTR_PT(451) OR ROM64_INSTR_PT(453)
     OR ROM64_INSTR_PT(454) OR ROM64_INSTR_PT(455)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(460) OR ROM64_INSTR_PT(463)
     OR ROM64_INSTR_PT(464) OR ROM64_INSTR_PT(466)
     OR ROM64_INSTR_PT(467) OR ROM64_INSTR_PT(468)
     OR ROM64_INSTR_PT(471) OR ROM64_INSTR_PT(472)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(474)
     OR ROM64_INSTR_PT(475) OR ROM64_INSTR_PT(483)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(491)
     OR ROM64_INSTR_PT(497) OR ROM64_INSTR_PT(498)
     OR ROM64_INSTR_PT(499) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(506) OR ROM64_INSTR_PT(508)
     OR ROM64_INSTR_PT(510) OR ROM64_INSTR_PT(514)
     OR ROM64_INSTR_PT(516) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(532) OR ROM64_INSTR_PT(538)
     OR ROM64_INSTR_PT(542) OR ROM64_INSTR_PT(546)
     OR ROM64_INSTR_PT(549) OR ROM64_INSTR_PT(551)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(559) OR ROM64_INSTR_PT(562)
     OR ROM64_INSTR_PT(566) OR ROM64_INSTR_PT(570)
     OR ROM64_INSTR_PT(571) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(581)
     OR ROM64_INSTR_PT(586) OR ROM64_INSTR_PT(589)
     OR ROM64_INSTR_PT(593) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(598)
     OR ROM64_INSTR_PT(601) OR ROM64_INSTR_PT(603)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(606)
     OR ROM64_INSTR_PT(611) OR ROM64_INSTR_PT(612)
     OR ROM64_INSTR_PT(613) OR ROM64_INSTR_PT(614)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(616)
     OR ROM64_INSTR_PT(617) OR ROM64_INSTR_PT(620)
     OR ROM64_INSTR_PT(626) OR ROM64_INSTR_PT(627)
     OR ROM64_INSTR_PT(628) OR ROM64_INSTR_PT(632)
     OR ROM64_INSTR_PT(635) OR ROM64_INSTR_PT(654)
     OR ROM64_INSTR_PT(659) OR ROM64_INSTR_PT(660)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(668)
     OR ROM64_INSTR_PT(675) OR ROM64_INSTR_PT(679)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(682)
     OR ROM64_INSTR_PT(687) OR ROM64_INSTR_PT(691)
     OR ROM64_INSTR_PT(703) OR ROM64_INSTR_PT(709)
     OR ROM64_INSTR_PT(711) OR ROM64_INSTR_PT(713)
     OR ROM64_INSTR_PT(717) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(728)
     OR ROM64_INSTR_PT(733) OR ROM64_INSTR_PT(735)
     OR ROM64_INSTR_PT(738) OR ROM64_INSTR_PT(741)
     OR ROM64_INSTR_PT(759) OR ROM64_INSTR_PT(766)
     OR ROM64_INSTR_PT(781) OR ROM64_INSTR_PT(791)
     OR ROM64_INSTR_PT(794) OR ROM64_INSTR_PT(797)
     OR ROM64_INSTR_PT(801) OR ROM64_INSTR_PT(808)
     OR ROM64_INSTR_PT(809) OR ROM64_INSTR_PT(811)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(822)
     OR ROM64_INSTR_PT(824) OR ROM64_INSTR_PT(846)
     OR ROM64_INSTR_PT(849) OR ROM64_INSTR_PT(852)
     OR ROM64_INSTR_PT(854) OR ROM64_INSTR_PT(855)
     OR ROM64_INSTR_PT(869) OR ROM64_INSTR_PT(872)
     OR ROM64_INSTR_PT(883) OR ROM64_INSTR_PT(886)
    );
MQQ894:TEMPLATE(3) <= 
    (ROM64_INSTR_PT(2) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(9)
     OR ROM64_INSTR_PT(10) OR ROM64_INSTR_PT(11)
     OR ROM64_INSTR_PT(14) OR ROM64_INSTR_PT(15)
     OR ROM64_INSTR_PT(17) OR ROM64_INSTR_PT(18)
     OR ROM64_INSTR_PT(20) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(25)
     OR ROM64_INSTR_PT(28) OR ROM64_INSTR_PT(29)
     OR ROM64_INSTR_PT(33) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(35) OR ROM64_INSTR_PT(36)
     OR ROM64_INSTR_PT(38) OR ROM64_INSTR_PT(39)
     OR ROM64_INSTR_PT(41) OR ROM64_INSTR_PT(42)
     OR ROM64_INSTR_PT(43) OR ROM64_INSTR_PT(45)
     OR ROM64_INSTR_PT(49) OR ROM64_INSTR_PT(52)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(56)
     OR ROM64_INSTR_PT(60) OR ROM64_INSTR_PT(61)
     OR ROM64_INSTR_PT(64) OR ROM64_INSTR_PT(66)
     OR ROM64_INSTR_PT(69) OR ROM64_INSTR_PT(70)
     OR ROM64_INSTR_PT(71) OR ROM64_INSTR_PT(73)
     OR ROM64_INSTR_PT(75) OR ROM64_INSTR_PT(76)
     OR ROM64_INSTR_PT(77) OR ROM64_INSTR_PT(78)
     OR ROM64_INSTR_PT(80) OR ROM64_INSTR_PT(82)
     OR ROM64_INSTR_PT(83) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(86) OR ROM64_INSTR_PT(89)
     OR ROM64_INSTR_PT(90) OR ROM64_INSTR_PT(92)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(95)
     OR ROM64_INSTR_PT(96) OR ROM64_INSTR_PT(97)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(99)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(102)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(106)
     OR ROM64_INSTR_PT(108) OR ROM64_INSTR_PT(109)
     OR ROM64_INSTR_PT(110) OR ROM64_INSTR_PT(113)
     OR ROM64_INSTR_PT(114) OR ROM64_INSTR_PT(115)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(124)
     OR ROM64_INSTR_PT(127) OR ROM64_INSTR_PT(133)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(140)
     OR ROM64_INSTR_PT(142) OR ROM64_INSTR_PT(144)
     OR ROM64_INSTR_PT(145) OR ROM64_INSTR_PT(146)
     OR ROM64_INSTR_PT(147) OR ROM64_INSTR_PT(148)
     OR ROM64_INSTR_PT(150) OR ROM64_INSTR_PT(151)
     OR ROM64_INSTR_PT(153) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(160) OR ROM64_INSTR_PT(161)
     OR ROM64_INSTR_PT(164) OR ROM64_INSTR_PT(166)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(169)
     OR ROM64_INSTR_PT(171) OR ROM64_INSTR_PT(172)
     OR ROM64_INSTR_PT(173) OR ROM64_INSTR_PT(174)
     OR ROM64_INSTR_PT(175) OR ROM64_INSTR_PT(177)
     OR ROM64_INSTR_PT(179) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(181) OR ROM64_INSTR_PT(182)
     OR ROM64_INSTR_PT(183) OR ROM64_INSTR_PT(184)
     OR ROM64_INSTR_PT(186) OR ROM64_INSTR_PT(187)
     OR ROM64_INSTR_PT(188) OR ROM64_INSTR_PT(191)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(199)
     OR ROM64_INSTR_PT(201) OR ROM64_INSTR_PT(202)
     OR ROM64_INSTR_PT(203) OR ROM64_INSTR_PT(205)
     OR ROM64_INSTR_PT(206) OR ROM64_INSTR_PT(207)
     OR ROM64_INSTR_PT(208) OR ROM64_INSTR_PT(209)
     OR ROM64_INSTR_PT(211) OR ROM64_INSTR_PT(215)
     OR ROM64_INSTR_PT(216) OR ROM64_INSTR_PT(217)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(219)
     OR ROM64_INSTR_PT(221) OR ROM64_INSTR_PT(222)
     OR ROM64_INSTR_PT(223) OR ROM64_INSTR_PT(225)
     OR ROM64_INSTR_PT(226) OR ROM64_INSTR_PT(228)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(231) OR ROM64_INSTR_PT(233)
     OR ROM64_INSTR_PT(238) OR ROM64_INSTR_PT(240)
     OR ROM64_INSTR_PT(242) OR ROM64_INSTR_PT(243)
     OR ROM64_INSTR_PT(245) OR ROM64_INSTR_PT(247)
     OR ROM64_INSTR_PT(249) OR ROM64_INSTR_PT(252)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(254)
     OR ROM64_INSTR_PT(257) OR ROM64_INSTR_PT(258)
     OR ROM64_INSTR_PT(259) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(265) OR ROM64_INSTR_PT(268)
     OR ROM64_INSTR_PT(269) OR ROM64_INSTR_PT(270)
     OR ROM64_INSTR_PT(271) OR ROM64_INSTR_PT(272)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(274)
     OR ROM64_INSTR_PT(275) OR ROM64_INSTR_PT(277)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(281)
     OR ROM64_INSTR_PT(282) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(287) OR ROM64_INSTR_PT(288)
     OR ROM64_INSTR_PT(290) OR ROM64_INSTR_PT(293)
     OR ROM64_INSTR_PT(294) OR ROM64_INSTR_PT(295)
     OR ROM64_INSTR_PT(298) OR ROM64_INSTR_PT(299)
     OR ROM64_INSTR_PT(302) OR ROM64_INSTR_PT(304)
     OR ROM64_INSTR_PT(305) OR ROM64_INSTR_PT(307)
     OR ROM64_INSTR_PT(309) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(313) OR ROM64_INSTR_PT(315)
     OR ROM64_INSTR_PT(319) OR ROM64_INSTR_PT(324)
     OR ROM64_INSTR_PT(325) OR ROM64_INSTR_PT(327)
     OR ROM64_INSTR_PT(331) OR ROM64_INSTR_PT(332)
     OR ROM64_INSTR_PT(334) OR ROM64_INSTR_PT(339)
     OR ROM64_INSTR_PT(340) OR ROM64_INSTR_PT(341)
     OR ROM64_INSTR_PT(342) OR ROM64_INSTR_PT(348)
     OR ROM64_INSTR_PT(350) OR ROM64_INSTR_PT(352)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(359)
     OR ROM64_INSTR_PT(361) OR ROM64_INSTR_PT(364)
     OR ROM64_INSTR_PT(365) OR ROM64_INSTR_PT(366)
     OR ROM64_INSTR_PT(369) OR ROM64_INSTR_PT(371)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(374)
     OR ROM64_INSTR_PT(375) OR ROM64_INSTR_PT(378)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(383) OR ROM64_INSTR_PT(384)
     OR ROM64_INSTR_PT(385) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(389) OR ROM64_INSTR_PT(391)
     OR ROM64_INSTR_PT(394) OR ROM64_INSTR_PT(395)
     OR ROM64_INSTR_PT(396) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(403)
     OR ROM64_INSTR_PT(404) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(406) OR ROM64_INSTR_PT(408)
     OR ROM64_INSTR_PT(409) OR ROM64_INSTR_PT(410)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(419) OR ROM64_INSTR_PT(420)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(424)
     OR ROM64_INSTR_PT(425) OR ROM64_INSTR_PT(426)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(428)
     OR ROM64_INSTR_PT(429) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(437) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(439) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(443)
     OR ROM64_INSTR_PT(445) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(448) OR ROM64_INSTR_PT(451)
     OR ROM64_INSTR_PT(453) OR ROM64_INSTR_PT(454)
     OR ROM64_INSTR_PT(455) OR ROM64_INSTR_PT(456)
     OR ROM64_INSTR_PT(457) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(460) OR ROM64_INSTR_PT(463)
     OR ROM64_INSTR_PT(464) OR ROM64_INSTR_PT(466)
     OR ROM64_INSTR_PT(467) OR ROM64_INSTR_PT(468)
     OR ROM64_INSTR_PT(470) OR ROM64_INSTR_PT(471)
     OR ROM64_INSTR_PT(472) OR ROM64_INSTR_PT(473)
     OR ROM64_INSTR_PT(474) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(478) OR ROM64_INSTR_PT(481)
     OR ROM64_INSTR_PT(482) OR ROM64_INSTR_PT(483)
     OR ROM64_INSTR_PT(484) OR ROM64_INSTR_PT(485)
     OR ROM64_INSTR_PT(488) OR ROM64_INSTR_PT(490)
     OR ROM64_INSTR_PT(491) OR ROM64_INSTR_PT(493)
     OR ROM64_INSTR_PT(495) OR ROM64_INSTR_PT(497)
     OR ROM64_INSTR_PT(498) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(505) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(508) OR ROM64_INSTR_PT(509)
     OR ROM64_INSTR_PT(510) OR ROM64_INSTR_PT(511)
     OR ROM64_INSTR_PT(516) OR ROM64_INSTR_PT(517)
     OR ROM64_INSTR_PT(519) OR ROM64_INSTR_PT(520)
     OR ROM64_INSTR_PT(521) OR ROM64_INSTR_PT(522)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(525)
     OR ROM64_INSTR_PT(532) OR ROM64_INSTR_PT(534)
     OR ROM64_INSTR_PT(538) OR ROM64_INSTR_PT(542)
     OR ROM64_INSTR_PT(546) OR ROM64_INSTR_PT(549)
     OR ROM64_INSTR_PT(551) OR ROM64_INSTR_PT(552)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(555) OR ROM64_INSTR_PT(558)
     OR ROM64_INSTR_PT(559) OR ROM64_INSTR_PT(562)
     OR ROM64_INSTR_PT(563) OR ROM64_INSTR_PT(564)
     OR ROM64_INSTR_PT(566) OR ROM64_INSTR_PT(569)
     OR ROM64_INSTR_PT(570) OR ROM64_INSTR_PT(571)
     OR ROM64_INSTR_PT(572) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(581)
     OR ROM64_INSTR_PT(582) OR ROM64_INSTR_PT(583)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(585)
     OR ROM64_INSTR_PT(586) OR ROM64_INSTR_PT(587)
     OR ROM64_INSTR_PT(588) OR ROM64_INSTR_PT(589)
     OR ROM64_INSTR_PT(590) OR ROM64_INSTR_PT(592)
     OR ROM64_INSTR_PT(595) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(598)
     OR ROM64_INSTR_PT(600) OR ROM64_INSTR_PT(601)
     OR ROM64_INSTR_PT(603) OR ROM64_INSTR_PT(604)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(610) OR ROM64_INSTR_PT(611)
     OR ROM64_INSTR_PT(612) OR ROM64_INSTR_PT(613)
     OR ROM64_INSTR_PT(614) OR ROM64_INSTR_PT(615)
     OR ROM64_INSTR_PT(616) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(620)
     OR ROM64_INSTR_PT(623) OR ROM64_INSTR_PT(626)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(629) OR ROM64_INSTR_PT(632)
     OR ROM64_INSTR_PT(633) OR ROM64_INSTR_PT(635)
     OR ROM64_INSTR_PT(636) OR ROM64_INSTR_PT(639)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(644)
     OR ROM64_INSTR_PT(654) OR ROM64_INSTR_PT(657)
     OR ROM64_INSTR_PT(659) OR ROM64_INSTR_PT(660)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(664)
     OR ROM64_INSTR_PT(666) OR ROM64_INSTR_PT(668)
     OR ROM64_INSTR_PT(675) OR ROM64_INSTR_PT(678)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(682)
     OR ROM64_INSTR_PT(691) OR ROM64_INSTR_PT(695)
     OR ROM64_INSTR_PT(703) OR ROM64_INSTR_PT(706)
     OR ROM64_INSTR_PT(709) OR ROM64_INSTR_PT(713)
     OR ROM64_INSTR_PT(717) OR ROM64_INSTR_PT(721)
     OR ROM64_INSTR_PT(722) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(728)
     OR ROM64_INSTR_PT(731) OR ROM64_INSTR_PT(733)
     OR ROM64_INSTR_PT(735) OR ROM64_INSTR_PT(736)
     OR ROM64_INSTR_PT(738) OR ROM64_INSTR_PT(744)
     OR ROM64_INSTR_PT(759) OR ROM64_INSTR_PT(761)
     OR ROM64_INSTR_PT(766) OR ROM64_INSTR_PT(769)
     OR ROM64_INSTR_PT(776) OR ROM64_INSTR_PT(781)
     OR ROM64_INSTR_PT(794) OR ROM64_INSTR_PT(797)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(809)
     OR ROM64_INSTR_PT(811) OR ROM64_INSTR_PT(813)
     OR ROM64_INSTR_PT(822) OR ROM64_INSTR_PT(824)
     OR ROM64_INSTR_PT(834) OR ROM64_INSTR_PT(846)
     OR ROM64_INSTR_PT(854) OR ROM64_INSTR_PT(855)
     OR ROM64_INSTR_PT(856) OR ROM64_INSTR_PT(858)
     OR ROM64_INSTR_PT(864) OR ROM64_INSTR_PT(869)
     OR ROM64_INSTR_PT(870) OR ROM64_INSTR_PT(883)
    );
MQQ895:TEMPLATE(4) <= 
    (ROM64_INSTR_PT(2) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(10)
     OR ROM64_INSTR_PT(14) OR ROM64_INSTR_PT(15)
     OR ROM64_INSTR_PT(18) OR ROM64_INSTR_PT(20)
     OR ROM64_INSTR_PT(25) OR ROM64_INSTR_PT(28)
     OR ROM64_INSTR_PT(29) OR ROM64_INSTR_PT(33)
     OR ROM64_INSTR_PT(35) OR ROM64_INSTR_PT(36)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(43)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(53)
     OR ROM64_INSTR_PT(56) OR ROM64_INSTR_PT(60)
     OR ROM64_INSTR_PT(65) OR ROM64_INSTR_PT(66)
     OR ROM64_INSTR_PT(69) OR ROM64_INSTR_PT(73)
     OR ROM64_INSTR_PT(74) OR ROM64_INSTR_PT(77)
     OR ROM64_INSTR_PT(78) OR ROM64_INSTR_PT(79)
     OR ROM64_INSTR_PT(80) OR ROM64_INSTR_PT(82)
     OR ROM64_INSTR_PT(84) OR ROM64_INSTR_PT(89)
     OR ROM64_INSTR_PT(92) OR ROM64_INSTR_PT(95)
     OR ROM64_INSTR_PT(96) OR ROM64_INSTR_PT(97)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(101)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(106)
     OR ROM64_INSTR_PT(108) OR ROM64_INSTR_PT(109)
     OR ROM64_INSTR_PT(110) OR ROM64_INSTR_PT(112)
     OR ROM64_INSTR_PT(114) OR ROM64_INSTR_PT(116)
     OR ROM64_INSTR_PT(119) OR ROM64_INSTR_PT(124)
     OR ROM64_INSTR_PT(129) OR ROM64_INSTR_PT(139)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(142)
     OR ROM64_INSTR_PT(143) OR ROM64_INSTR_PT(145)
     OR ROM64_INSTR_PT(146) OR ROM64_INSTR_PT(147)
     OR ROM64_INSTR_PT(150) OR ROM64_INSTR_PT(151)
     OR ROM64_INSTR_PT(153) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(158) OR ROM64_INSTR_PT(160)
     OR ROM64_INSTR_PT(161) OR ROM64_INSTR_PT(166)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(172)
     OR ROM64_INSTR_PT(173) OR ROM64_INSTR_PT(174)
     OR ROM64_INSTR_PT(175) OR ROM64_INSTR_PT(176)
     OR ROM64_INSTR_PT(177) OR ROM64_INSTR_PT(179)
     OR ROM64_INSTR_PT(181) OR ROM64_INSTR_PT(182)
     OR ROM64_INSTR_PT(183) OR ROM64_INSTR_PT(184)
     OR ROM64_INSTR_PT(187) OR ROM64_INSTR_PT(188)
     OR ROM64_INSTR_PT(191) OR ROM64_INSTR_PT(193)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(202)
     OR ROM64_INSTR_PT(203) OR ROM64_INSTR_PT(205)
     OR ROM64_INSTR_PT(206) OR ROM64_INSTR_PT(207)
     OR ROM64_INSTR_PT(208) OR ROM64_INSTR_PT(209)
     OR ROM64_INSTR_PT(211) OR ROM64_INSTR_PT(216)
     OR ROM64_INSTR_PT(219) OR ROM64_INSTR_PT(221)
     OR ROM64_INSTR_PT(225) OR ROM64_INSTR_PT(228)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(231) OR ROM64_INSTR_PT(233)
     OR ROM64_INSTR_PT(237) OR ROM64_INSTR_PT(240)
     OR ROM64_INSTR_PT(242) OR ROM64_INSTR_PT(243)
     OR ROM64_INSTR_PT(247) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(254) OR ROM64_INSTR_PT(257)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(259)
     OR ROM64_INSTR_PT(260) OR ROM64_INSTR_PT(261)
     OR ROM64_INSTR_PT(265) OR ROM64_INSTR_PT(269)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(274)
     OR ROM64_INSTR_PT(277) OR ROM64_INSTR_PT(281)
     OR ROM64_INSTR_PT(284) OR ROM64_INSTR_PT(288)
     OR ROM64_INSTR_PT(290) OR ROM64_INSTR_PT(292)
     OR ROM64_INSTR_PT(294) OR ROM64_INSTR_PT(295)
     OR ROM64_INSTR_PT(304) OR ROM64_INSTR_PT(307)
     OR ROM64_INSTR_PT(309) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(313) OR ROM64_INSTR_PT(319)
     OR ROM64_INSTR_PT(320) OR ROM64_INSTR_PT(324)
     OR ROM64_INSTR_PT(325) OR ROM64_INSTR_PT(327)
     OR ROM64_INSTR_PT(332) OR ROM64_INSTR_PT(334)
     OR ROM64_INSTR_PT(339) OR ROM64_INSTR_PT(340)
     OR ROM64_INSTR_PT(341) OR ROM64_INSTR_PT(342)
     OR ROM64_INSTR_PT(348) OR ROM64_INSTR_PT(350)
     OR ROM64_INSTR_PT(352) OR ROM64_INSTR_PT(353)
     OR ROM64_INSTR_PT(358) OR ROM64_INSTR_PT(359)
     OR ROM64_INSTR_PT(360) OR ROM64_INSTR_PT(361)
     OR ROM64_INSTR_PT(362) OR ROM64_INSTR_PT(365)
     OR ROM64_INSTR_PT(366) OR ROM64_INSTR_PT(368)
     OR ROM64_INSTR_PT(369) OR ROM64_INSTR_PT(371)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(374)
     OR ROM64_INSTR_PT(377) OR ROM64_INSTR_PT(378)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(389) OR ROM64_INSTR_PT(392)
     OR ROM64_INSTR_PT(394) OR ROM64_INSTR_PT(395)
     OR ROM64_INSTR_PT(396) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(402) OR ROM64_INSTR_PT(403)
     OR ROM64_INSTR_PT(405) OR ROM64_INSTR_PT(406)
     OR ROM64_INSTR_PT(408) OR ROM64_INSTR_PT(409)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(419) OR ROM64_INSTR_PT(420)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(425)
     OR ROM64_INSTR_PT(426) OR ROM64_INSTR_PT(428)
     OR ROM64_INSTR_PT(429) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(438) OR ROM64_INSTR_PT(439)
     OR ROM64_INSTR_PT(440) OR ROM64_INSTR_PT(443)
     OR ROM64_INSTR_PT(445) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(448) OR ROM64_INSTR_PT(451)
     OR ROM64_INSTR_PT(453) OR ROM64_INSTR_PT(454)
     OR ROM64_INSTR_PT(455) OR ROM64_INSTR_PT(456)
     OR ROM64_INSTR_PT(458) OR ROM64_INSTR_PT(460)
     OR ROM64_INSTR_PT(463) OR ROM64_INSTR_PT(464)
     OR ROM64_INSTR_PT(466) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(468) OR ROM64_INSTR_PT(470)
     OR ROM64_INSTR_PT(471) OR ROM64_INSTR_PT(472)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(474)
     OR ROM64_INSTR_PT(475) OR ROM64_INSTR_PT(477)
     OR ROM64_INSTR_PT(483) OR ROM64_INSTR_PT(490)
     OR ROM64_INSTR_PT(491) OR ROM64_INSTR_PT(497)
     OR ROM64_INSTR_PT(498) OR ROM64_INSTR_PT(499)
     OR ROM64_INSTR_PT(503) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(508) OR ROM64_INSTR_PT(510)
     OR ROM64_INSTR_PT(516) OR ROM64_INSTR_PT(517)
     OR ROM64_INSTR_PT(519) OR ROM64_INSTR_PT(520)
     OR ROM64_INSTR_PT(527) OR ROM64_INSTR_PT(532)
     OR ROM64_INSTR_PT(538) OR ROM64_INSTR_PT(542)
     OR ROM64_INSTR_PT(546) OR ROM64_INSTR_PT(549)
     OR ROM64_INSTR_PT(551) OR ROM64_INSTR_PT(553)
     OR ROM64_INSTR_PT(554) OR ROM64_INSTR_PT(557)
     OR ROM64_INSTR_PT(559) OR ROM64_INSTR_PT(562)
     OR ROM64_INSTR_PT(564) OR ROM64_INSTR_PT(566)
     OR ROM64_INSTR_PT(570) OR ROM64_INSTR_PT(571)
     OR ROM64_INSTR_PT(572) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(581)
     OR ROM64_INSTR_PT(586) OR ROM64_INSTR_PT(589)
     OR ROM64_INSTR_PT(590) OR ROM64_INSTR_PT(593)
     OR ROM64_INSTR_PT(596) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(598) OR ROM64_INSTR_PT(601)
     OR ROM64_INSTR_PT(602) OR ROM64_INSTR_PT(603)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(606)
     OR ROM64_INSTR_PT(610) OR ROM64_INSTR_PT(611)
     OR ROM64_INSTR_PT(612) OR ROM64_INSTR_PT(613)
     OR ROM64_INSTR_PT(614) OR ROM64_INSTR_PT(615)
     OR ROM64_INSTR_PT(616) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(620) OR ROM64_INSTR_PT(626)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(632) OR ROM64_INSTR_PT(635)
     OR ROM64_INSTR_PT(636) OR ROM64_INSTR_PT(641)
     OR ROM64_INSTR_PT(653) OR ROM64_INSTR_PT(654)
     OR ROM64_INSTR_PT(659) OR ROM64_INSTR_PT(660)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(664)
     OR ROM64_INSTR_PT(668) OR ROM64_INSTR_PT(675)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(682)
     OR ROM64_INSTR_PT(685) OR ROM64_INSTR_PT(691)
     OR ROM64_INSTR_PT(694) OR ROM64_INSTR_PT(695)
     OR ROM64_INSTR_PT(702) OR ROM64_INSTR_PT(703)
     OR ROM64_INSTR_PT(706) OR ROM64_INSTR_PT(709)
     OR ROM64_INSTR_PT(713) OR ROM64_INSTR_PT(716)
     OR ROM64_INSTR_PT(717) OR ROM64_INSTR_PT(721)
     OR ROM64_INSTR_PT(723) OR ROM64_INSTR_PT(724)
     OR ROM64_INSTR_PT(728) OR ROM64_INSTR_PT(733)
     OR ROM64_INSTR_PT(735) OR ROM64_INSTR_PT(736)
     OR ROM64_INSTR_PT(738) OR ROM64_INSTR_PT(741)
     OR ROM64_INSTR_PT(759) OR ROM64_INSTR_PT(766)
     OR ROM64_INSTR_PT(770) OR ROM64_INSTR_PT(781)
     OR ROM64_INSTR_PT(794) OR ROM64_INSTR_PT(797)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(801)
     OR ROM64_INSTR_PT(808) OR ROM64_INSTR_PT(809)
     OR ROM64_INSTR_PT(811) OR ROM64_INSTR_PT(813)
     OR ROM64_INSTR_PT(822) OR ROM64_INSTR_PT(824)
     OR ROM64_INSTR_PT(832) OR ROM64_INSTR_PT(834)
     OR ROM64_INSTR_PT(846) OR ROM64_INSTR_PT(849)
     OR ROM64_INSTR_PT(852) OR ROM64_INSTR_PT(854)
     OR ROM64_INSTR_PT(855) OR ROM64_INSTR_PT(858)
     OR ROM64_INSTR_PT(869) OR ROM64_INSTR_PT(873)
     OR ROM64_INSTR_PT(883));
MQQ896:TEMPLATE(5) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(6)
     OR ROM64_INSTR_PT(7) OR ROM64_INSTR_PT(8)
     OR ROM64_INSTR_PT(11) OR ROM64_INSTR_PT(14)
     OR ROM64_INSTR_PT(15) OR ROM64_INSTR_PT(18)
     OR ROM64_INSTR_PT(21) OR ROM64_INSTR_PT(35)
     OR ROM64_INSTR_PT(38) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(45)
     OR ROM64_INSTR_PT(49) OR ROM64_INSTR_PT(51)
     OR ROM64_INSTR_PT(52) OR ROM64_INSTR_PT(53)
     OR ROM64_INSTR_PT(56) OR ROM64_INSTR_PT(57)
     OR ROM64_INSTR_PT(61) OR ROM64_INSTR_PT(64)
     OR ROM64_INSTR_PT(68) OR ROM64_INSTR_PT(69)
     OR ROM64_INSTR_PT(70) OR ROM64_INSTR_PT(73)
     OR ROM64_INSTR_PT(82) OR ROM64_INSTR_PT(83)
     OR ROM64_INSTR_PT(84) OR ROM64_INSTR_PT(86)
     OR ROM64_INSTR_PT(90) OR ROM64_INSTR_PT(93)
     OR ROM64_INSTR_PT(95) OR ROM64_INSTR_PT(100)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(102)
     OR ROM64_INSTR_PT(105) OR ROM64_INSTR_PT(108)
     OR ROM64_INSTR_PT(109) OR ROM64_INSTR_PT(115)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(124)
     OR ROM64_INSTR_PT(128) OR ROM64_INSTR_PT(132)
     OR ROM64_INSTR_PT(133) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(143)
     OR ROM64_INSTR_PT(144) OR ROM64_INSTR_PT(145)
     OR ROM64_INSTR_PT(153) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(157) OR ROM64_INSTR_PT(158)
     OR ROM64_INSTR_PT(162) OR ROM64_INSTR_PT(164)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(169)
     OR ROM64_INSTR_PT(170) OR ROM64_INSTR_PT(177)
     OR ROM64_INSTR_PT(180) OR ROM64_INSTR_PT(181)
     OR ROM64_INSTR_PT(183) OR ROM64_INSTR_PT(185)
     OR ROM64_INSTR_PT(186) OR ROM64_INSTR_PT(194)
     OR ROM64_INSTR_PT(196) OR ROM64_INSTR_PT(201)
     OR ROM64_INSTR_PT(203) OR ROM64_INSTR_PT(204)
     OR ROM64_INSTR_PT(205) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(211) OR ROM64_INSTR_PT(215)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(219)
     OR ROM64_INSTR_PT(223) OR ROM64_INSTR_PT(226)
     OR ROM64_INSTR_PT(233) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(241) OR ROM64_INSTR_PT(243)
     OR ROM64_INSTR_PT(244) OR ROM64_INSTR_PT(245)
     OR ROM64_INSTR_PT(249) OR ROM64_INSTR_PT(254)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(263) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(265) OR ROM64_INSTR_PT(268)
     OR ROM64_INSTR_PT(269) OR ROM64_INSTR_PT(270)
     OR ROM64_INSTR_PT(272) OR ROM64_INSTR_PT(276)
     OR ROM64_INSTR_PT(278) OR ROM64_INSTR_PT(280)
     OR ROM64_INSTR_PT(282) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(285) OR ROM64_INSTR_PT(287)
     OR ROM64_INSTR_PT(290) OR ROM64_INSTR_PT(293)
     OR ROM64_INSTR_PT(294) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(302) OR ROM64_INSTR_PT(305)
     OR ROM64_INSTR_PT(308) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(312) OR ROM64_INSTR_PT(319)
     OR ROM64_INSTR_PT(325) OR ROM64_INSTR_PT(339)
     OR ROM64_INSTR_PT(348) OR ROM64_INSTR_PT(350)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(355)
     OR ROM64_INSTR_PT(358) OR ROM64_INSTR_PT(364)
     OR ROM64_INSTR_PT(366) OR ROM64_INSTR_PT(367)
     OR ROM64_INSTR_PT(370) OR ROM64_INSTR_PT(372)
     OR ROM64_INSTR_PT(375) OR ROM64_INSTR_PT(378)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(383)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(385)
     OR ROM64_INSTR_PT(391) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(399) OR ROM64_INSTR_PT(403)
     OR ROM64_INSTR_PT(405) OR ROM64_INSTR_PT(409)
     OR ROM64_INSTR_PT(410) OR ROM64_INSTR_PT(413)
     OR ROM64_INSTR_PT(416) OR ROM64_INSTR_PT(417)
     OR ROM64_INSTR_PT(418) OR ROM64_INSTR_PT(419)
     OR ROM64_INSTR_PT(425) OR ROM64_INSTR_PT(426)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(428)
     OR ROM64_INSTR_PT(429) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(432) OR ROM64_INSTR_PT(433)
     OR ROM64_INSTR_PT(435) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(439) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(443)
     OR ROM64_INSTR_PT(445) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(451) OR ROM64_INSTR_PT(453)
     OR ROM64_INSTR_PT(454) OR ROM64_INSTR_PT(455)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(457)
     OR ROM64_INSTR_PT(460) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(478) OR ROM64_INSTR_PT(481)
     OR ROM64_INSTR_PT(482) OR ROM64_INSTR_PT(484)
     OR ROM64_INSTR_PT(485) OR ROM64_INSTR_PT(488)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(493)
     OR ROM64_INSTR_PT(495) OR ROM64_INSTR_PT(496)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(510) OR ROM64_INSTR_PT(512)
     OR ROM64_INSTR_PT(514) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(522) OR ROM64_INSTR_PT(523)
     OR ROM64_INSTR_PT(525) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(531) OR ROM64_INSTR_PT(532)
     OR ROM64_INSTR_PT(534) OR ROM64_INSTR_PT(539)
     OR ROM64_INSTR_PT(542) OR ROM64_INSTR_PT(546)
     OR ROM64_INSTR_PT(552) OR ROM64_INSTR_PT(553)
     OR ROM64_INSTR_PT(554) OR ROM64_INSTR_PT(555)
     OR ROM64_INSTR_PT(557) OR ROM64_INSTR_PT(559)
     OR ROM64_INSTR_PT(563) OR ROM64_INSTR_PT(564)
     OR ROM64_INSTR_PT(566) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(570) OR ROM64_INSTR_PT(571)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(577)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(581)
     OR ROM64_INSTR_PT(582) OR ROM64_INSTR_PT(583)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(585)
     OR ROM64_INSTR_PT(586) OR ROM64_INSTR_PT(587)
     OR ROM64_INSTR_PT(589) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(592) OR ROM64_INSTR_PT(604)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(607)
     OR ROM64_INSTR_PT(608) OR ROM64_INSTR_PT(611)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(616)
     OR ROM64_INSTR_PT(619) OR ROM64_INSTR_PT(625)
     OR ROM64_INSTR_PT(626) OR ROM64_INSTR_PT(627)
     OR ROM64_INSTR_PT(629) OR ROM64_INSTR_PT(633)
     OR ROM64_INSTR_PT(636) OR ROM64_INSTR_PT(639)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(643)
     OR ROM64_INSTR_PT(655) OR ROM64_INSTR_PT(660)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(664)
     OR ROM64_INSTR_PT(666) OR ROM64_INSTR_PT(678)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(695)
     OR ROM64_INSTR_PT(698) OR ROM64_INSTR_PT(702)
     OR ROM64_INSTR_PT(713) OR ROM64_INSTR_PT(716)
     OR ROM64_INSTR_PT(721) OR ROM64_INSTR_PT(722)
     OR ROM64_INSTR_PT(731) OR ROM64_INSTR_PT(736)
     OR ROM64_INSTR_PT(753) OR ROM64_INSTR_PT(761)
     OR ROM64_INSTR_PT(769) OR ROM64_INSTR_PT(770)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(811)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(823)
     OR ROM64_INSTR_PT(824) OR ROM64_INSTR_PT(832)
     OR ROM64_INSTR_PT(834) OR ROM64_INSTR_PT(846)
     OR ROM64_INSTR_PT(854) OR ROM64_INSTR_PT(855)
     OR ROM64_INSTR_PT(856) OR ROM64_INSTR_PT(858)
     OR ROM64_INSTR_PT(864) OR ROM64_INSTR_PT(870)
     OR ROM64_INSTR_PT(873));
MQQ897:TEMPLATE(6) <= 
    ('0');
MQQ898:TEMPLATE(7) <= 
    ('0');
MQQ899:TEMPLATE(8) <= 
    ('0');
MQQ900:TEMPLATE(9) <= 
    (ROM64_INSTR_PT(7) OR ROM64_INSTR_PT(9)
     OR ROM64_INSTR_PT(11) OR ROM64_INSTR_PT(13)
     OR ROM64_INSTR_PT(15) OR ROM64_INSTR_PT(22)
     OR ROM64_INSTR_PT(25) OR ROM64_INSTR_PT(29)
     OR ROM64_INSTR_PT(36) OR ROM64_INSTR_PT(38)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(45)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(55)
     OR ROM64_INSTR_PT(56) OR ROM64_INSTR_PT(58)
     OR ROM64_INSTR_PT(61) OR ROM64_INSTR_PT(70)
     OR ROM64_INSTR_PT(71) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(86) OR ROM64_INSTR_PT(90)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(97)
     OR ROM64_INSTR_PT(100) OR ROM64_INSTR_PT(102)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(105)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(119)
     OR ROM64_INSTR_PT(124) OR ROM64_INSTR_PT(132)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(143) OR ROM64_INSTR_PT(144)
     OR ROM64_INSTR_PT(148) OR ROM64_INSTR_PT(154)
     OR ROM64_INSTR_PT(155) OR ROM64_INSTR_PT(160)
     OR ROM64_INSTR_PT(172) OR ROM64_INSTR_PT(174)
     OR ROM64_INSTR_PT(176) OR ROM64_INSTR_PT(177)
     OR ROM64_INSTR_PT(179) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(181) OR ROM64_INSTR_PT(183)
     OR ROM64_INSTR_PT(186) OR ROM64_INSTR_PT(193)
     OR ROM64_INSTR_PT(201) OR ROM64_INSTR_PT(208)
     OR ROM64_INSTR_PT(213) OR ROM64_INSTR_PT(215)
     OR ROM64_INSTR_PT(216) OR ROM64_INSTR_PT(221)
     OR ROM64_INSTR_PT(222) OR ROM64_INSTR_PT(225)
     OR ROM64_INSTR_PT(226) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(240) OR ROM64_INSTR_PT(242)
     OR ROM64_INSTR_PT(243) OR ROM64_INSTR_PT(245)
     OR ROM64_INSTR_PT(249) OR ROM64_INSTR_PT(259)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(262)
     OR ROM64_INSTR_PT(263) OR ROM64_INSTR_PT(265)
     OR ROM64_INSTR_PT(270) OR ROM64_INSTR_PT(274)
     OR ROM64_INSTR_PT(275) OR ROM64_INSTR_PT(276)
     OR ROM64_INSTR_PT(277) OR ROM64_INSTR_PT(282)
     OR ROM64_INSTR_PT(284) OR ROM64_INSTR_PT(285)
     OR ROM64_INSTR_PT(286) OR ROM64_INSTR_PT(292)
     OR ROM64_INSTR_PT(293) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(299) OR ROM64_INSTR_PT(302)
     OR ROM64_INSTR_PT(305) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(315) OR ROM64_INSTR_PT(319)
     OR ROM64_INSTR_PT(320) OR ROM64_INSTR_PT(322)
     OR ROM64_INSTR_PT(341) OR ROM64_INSTR_PT(349)
     OR ROM64_INSTR_PT(355) OR ROM64_INSTR_PT(359)
     OR ROM64_INSTR_PT(362) OR ROM64_INSTR_PT(365)
     OR ROM64_INSTR_PT(366) OR ROM64_INSTR_PT(369)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(379)
     OR ROM64_INSTR_PT(382) OR ROM64_INSTR_PT(383)
     OR ROM64_INSTR_PT(385) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(389) OR ROM64_INSTR_PT(392)
     OR ROM64_INSTR_PT(394) OR ROM64_INSTR_PT(395)
     OR ROM64_INSTR_PT(396) OR ROM64_INSTR_PT(402)
     OR ROM64_INSTR_PT(403) OR ROM64_INSTR_PT(404)
     OR ROM64_INSTR_PT(405) OR ROM64_INSTR_PT(410)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(415)
     OR ROM64_INSTR_PT(418) OR ROM64_INSTR_PT(425)
     OR ROM64_INSTR_PT(426) OR ROM64_INSTR_PT(429)
     OR ROM64_INSTR_PT(434) OR ROM64_INSTR_PT(435)
     OR ROM64_INSTR_PT(437) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(440) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(451)
     OR ROM64_INSTR_PT(453) OR ROM64_INSTR_PT(456)
     OR ROM64_INSTR_PT(457) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(470) OR ROM64_INSTR_PT(473)
     OR ROM64_INSTR_PT(474) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(478) OR ROM64_INSTR_PT(482)
     OR ROM64_INSTR_PT(485) OR ROM64_INSTR_PT(491)
     OR ROM64_INSTR_PT(493) OR ROM64_INSTR_PT(495)
     OR ROM64_INSTR_PT(498) OR ROM64_INSTR_PT(499)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(505)
     OR ROM64_INSTR_PT(507) OR ROM64_INSTR_PT(509)
     OR ROM64_INSTR_PT(517) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(520) OR ROM64_INSTR_PT(521)
     OR ROM64_INSTR_PT(522) OR ROM64_INSTR_PT(532)
     OR ROM64_INSTR_PT(534) OR ROM64_INSTR_PT(535)
     OR ROM64_INSTR_PT(544) OR ROM64_INSTR_PT(546)
     OR ROM64_INSTR_PT(549) OR ROM64_INSTR_PT(552)
     OR ROM64_INSTR_PT(555) OR ROM64_INSTR_PT(558)
     OR ROM64_INSTR_PT(559) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(569) OR ROM64_INSTR_PT(571)
     OR ROM64_INSTR_PT(572) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(590)
     OR ROM64_INSTR_PT(591) OR ROM64_INSTR_PT(592)
     OR ROM64_INSTR_PT(593) OR ROM64_INSTR_PT(595)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(610) OR ROM64_INSTR_PT(612)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(623)
     OR ROM64_INSTR_PT(628) OR ROM64_INSTR_PT(633)
     OR ROM64_INSTR_PT(639) OR ROM64_INSTR_PT(645)
     OR ROM64_INSTR_PT(646) OR ROM64_INSTR_PT(653)
     OR ROM64_INSTR_PT(659) OR ROM64_INSTR_PT(663)
     OR ROM64_INSTR_PT(666) OR ROM64_INSTR_PT(678)
     OR ROM64_INSTR_PT(691) OR ROM64_INSTR_PT(693)
     OR ROM64_INSTR_PT(703) OR ROM64_INSTR_PT(705)
     OR ROM64_INSTR_PT(741) OR ROM64_INSTR_PT(753)
     OR ROM64_INSTR_PT(797) OR ROM64_INSTR_PT(846)
    );
MQQ901:TEMPLATE(10) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(6)
     OR ROM64_INSTR_PT(7) OR ROM64_INSTR_PT(14)
     OR ROM64_INSTR_PT(15) OR ROM64_INSTR_PT(17)
     OR ROM64_INSTR_PT(20) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(45)
     OR ROM64_INSTR_PT(51) OR ROM64_INSTR_PT(52)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(57)
     OR ROM64_INSTR_PT(73) OR ROM64_INSTR_PT(74)
     OR ROM64_INSTR_PT(75) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(99)
     OR ROM64_INSTR_PT(112) OR ROM64_INSTR_PT(113)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(122) OR ROM64_INSTR_PT(125)
     OR ROM64_INSTR_PT(127) OR ROM64_INSTR_PT(128)
     OR ROM64_INSTR_PT(129) OR ROM64_INSTR_PT(132)
     OR ROM64_INSTR_PT(139) OR ROM64_INSTR_PT(140)
     OR ROM64_INSTR_PT(143) OR ROM64_INSTR_PT(153)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(169)
     OR ROM64_INSTR_PT(171) OR ROM64_INSTR_PT(173)
     OR ROM64_INSTR_PT(174) OR ROM64_INSTR_PT(181)
     OR ROM64_INSTR_PT(183) OR ROM64_INSTR_PT(184)
     OR ROM64_INSTR_PT(185) OR ROM64_INSTR_PT(191)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(199)
     OR ROM64_INSTR_PT(202) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(204) OR ROM64_INSTR_PT(213)
     OR ROM64_INSTR_PT(217) OR ROM64_INSTR_PT(219)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(237) OR ROM64_INSTR_PT(240)
     OR ROM64_INSTR_PT(241) OR ROM64_INSTR_PT(252)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(258)
     OR ROM64_INSTR_PT(260) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(271)
     OR ROM64_INSTR_PT(272) OR ROM64_INSTR_PT(273)
     OR ROM64_INSTR_PT(276) OR ROM64_INSTR_PT(278)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(331)
     OR ROM64_INSTR_PT(339) OR ROM64_INSTR_PT(361)
     OR ROM64_INSTR_PT(364) OR ROM64_INSTR_PT(366)
     OR ROM64_INSTR_PT(367) OR ROM64_INSTR_PT(368)
     OR ROM64_INSTR_PT(374) OR ROM64_INSTR_PT(375)
     OR ROM64_INSTR_PT(377) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(391)
     OR ROM64_INSTR_PT(396) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(403) OR ROM64_INSTR_PT(406)
     OR ROM64_INSTR_PT(408) OR ROM64_INSTR_PT(420)
     OR ROM64_INSTR_PT(424) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(442) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(448) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(472) OR ROM64_INSTR_PT(477)
     OR ROM64_INSTR_PT(480) OR ROM64_INSTR_PT(481)
     OR ROM64_INSTR_PT(483) OR ROM64_INSTR_PT(491)
     OR ROM64_INSTR_PT(503) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(507) OR ROM64_INSTR_PT(508)
     OR ROM64_INSTR_PT(511) OR ROM64_INSTR_PT(512)
     OR ROM64_INSTR_PT(519) OR ROM64_INSTR_PT(525)
     OR ROM64_INSTR_PT(527) OR ROM64_INSTR_PT(531)
     OR ROM64_INSTR_PT(532) OR ROM64_INSTR_PT(538)
     OR ROM64_INSTR_PT(539) OR ROM64_INSTR_PT(545)
     OR ROM64_INSTR_PT(548) OR ROM64_INSTR_PT(553)
     OR ROM64_INSTR_PT(554) OR ROM64_INSTR_PT(557)
     OR ROM64_INSTR_PT(562) OR ROM64_INSTR_PT(563)
     OR ROM64_INSTR_PT(571) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(583) OR ROM64_INSTR_PT(588)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(599)
     OR ROM64_INSTR_PT(600) OR ROM64_INSTR_PT(602)
     OR ROM64_INSTR_PT(603) OR ROM64_INSTR_PT(609)
     OR ROM64_INSTR_PT(614) OR ROM64_INSTR_PT(619)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(629)
     OR ROM64_INSTR_PT(632) OR ROM64_INSTR_PT(636)
     OR ROM64_INSTR_PT(637) OR ROM64_INSTR_PT(641)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(644)
     OR ROM64_INSTR_PT(655) OR ROM64_INSTR_PT(682)
     OR ROM64_INSTR_PT(685) OR ROM64_INSTR_PT(691)
     OR ROM64_INSTR_PT(713) OR ROM64_INSTR_PT(717)
     OR ROM64_INSTR_PT(721) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(728)
     OR ROM64_INSTR_PT(733) OR ROM64_INSTR_PT(735)
     OR ROM64_INSTR_PT(736) OR ROM64_INSTR_PT(738)
     OR ROM64_INSTR_PT(739) OR ROM64_INSTR_PT(761)
     OR ROM64_INSTR_PT(770) OR ROM64_INSTR_PT(824)
     OR ROM64_INSTR_PT(858) OR ROM64_INSTR_PT(873)
    );
MQQ902:TEMPLATE(11) <= 
    ('0');
MQQ903:TEMPLATE(12) <= 
    ('0');
MQQ904:TEMPLATE(13) <= 
    ('0');
MQQ905:TEMPLATE(14) <= 
    (ROM64_INSTR_PT(7) OR ROM64_INSTR_PT(11)
     OR ROM64_INSTR_PT(13) OR ROM64_INSTR_PT(15)
     OR ROM64_INSTR_PT(17) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(25) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(36) OR ROM64_INSTR_PT(38)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(52)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(55)
     OR ROM64_INSTR_PT(56) OR ROM64_INSTR_PT(61)
     OR ROM64_INSTR_PT(64) OR ROM64_INSTR_PT(70)
     OR ROM64_INSTR_PT(73) OR ROM64_INSTR_PT(75)
     OR ROM64_INSTR_PT(77) OR ROM64_INSTR_PT(80)
     OR ROM64_INSTR_PT(84) OR ROM64_INSTR_PT(86)
     OR ROM64_INSTR_PT(89) OR ROM64_INSTR_PT(90)
     OR ROM64_INSTR_PT(92) OR ROM64_INSTR_PT(93)
     OR ROM64_INSTR_PT(96) OR ROM64_INSTR_PT(97)
     OR ROM64_INSTR_PT(99) OR ROM64_INSTR_PT(102)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(106)
     OR ROM64_INSTR_PT(110) OR ROM64_INSTR_PT(113)
     OR ROM64_INSTR_PT(114) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(125)
     OR ROM64_INSTR_PT(127) OR ROM64_INSTR_PT(128)
     OR ROM64_INSTR_PT(132) OR ROM64_INSTR_PT(139)
     OR ROM64_INSTR_PT(144) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(169) OR ROM64_INSTR_PT(171)
     OR ROM64_INSTR_PT(172) OR ROM64_INSTR_PT(174)
     OR ROM64_INSTR_PT(180) OR ROM64_INSTR_PT(181)
     OR ROM64_INSTR_PT(184) OR ROM64_INSTR_PT(186)
     OR ROM64_INSTR_PT(196) OR ROM64_INSTR_PT(199)
     OR ROM64_INSTR_PT(201) OR ROM64_INSTR_PT(202)
     OR ROM64_INSTR_PT(208) OR ROM64_INSTR_PT(213)
     OR ROM64_INSTR_PT(215) OR ROM64_INSTR_PT(216)
     OR ROM64_INSTR_PT(217) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(226) OR ROM64_INSTR_PT(229)
     OR ROM64_INSTR_PT(230) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(240) OR ROM64_INSTR_PT(252)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(270)
     OR ROM64_INSTR_PT(271) OR ROM64_INSTR_PT(272)
     OR ROM64_INSTR_PT(274) OR ROM64_INSTR_PT(275)
     OR ROM64_INSTR_PT(276) OR ROM64_INSTR_PT(277)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(282)
     OR ROM64_INSTR_PT(286) OR ROM64_INSTR_PT(287)
     OR ROM64_INSTR_PT(293) OR ROM64_INSTR_PT(294)
     OR ROM64_INSTR_PT(298) OR ROM64_INSTR_PT(302)
     OR ROM64_INSTR_PT(305) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(315) OR ROM64_INSTR_PT(322)
     OR ROM64_INSTR_PT(331) OR ROM64_INSTR_PT(349)
     OR ROM64_INSTR_PT(364) OR ROM64_INSTR_PT(365)
     OR ROM64_INSTR_PT(366) OR ROM64_INSTR_PT(369)
     OR ROM64_INSTR_PT(371) OR ROM64_INSTR_PT(372)
     OR ROM64_INSTR_PT(375) OR ROM64_INSTR_PT(377)
     OR ROM64_INSTR_PT(383) OR ROM64_INSTR_PT(385)
     OR ROM64_INSTR_PT(388) OR ROM64_INSTR_PT(391)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(396)
     OR ROM64_INSTR_PT(397) OR ROM64_INSTR_PT(403)
     OR ROM64_INSTR_PT(404) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(410) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(420)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(424)
     OR ROM64_INSTR_PT(426) OR ROM64_INSTR_PT(427)
     OR ROM64_INSTR_PT(434) OR ROM64_INSTR_PT(437)
     OR ROM64_INSTR_PT(440) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(457)
     OR ROM64_INSTR_PT(466) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(478) OR ROM64_INSTR_PT(482)
     OR ROM64_INSTR_PT(483) OR ROM64_INSTR_PT(484)
     OR ROM64_INSTR_PT(485) OR ROM64_INSTR_PT(488)
     OR ROM64_INSTR_PT(493) OR ROM64_INSTR_PT(495)
     OR ROM64_INSTR_PT(498) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(505) OR ROM64_INSTR_PT(511)
     OR ROM64_INSTR_PT(517) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(520) OR ROM64_INSTR_PT(521)
     OR ROM64_INSTR_PT(522) OR ROM64_INSTR_PT(523)
     OR ROM64_INSTR_PT(525) OR ROM64_INSTR_PT(532)
     OR ROM64_INSTR_PT(534) OR ROM64_INSTR_PT(535)
     OR ROM64_INSTR_PT(537) OR ROM64_INSTR_PT(539)
     OR ROM64_INSTR_PT(542) OR ROM64_INSTR_PT(544)
     OR ROM64_INSTR_PT(545) OR ROM64_INSTR_PT(548)
     OR ROM64_INSTR_PT(549) OR ROM64_INSTR_PT(552)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(555) OR ROM64_INSTR_PT(558)
     OR ROM64_INSTR_PT(568) OR ROM64_INSTR_PT(569)
     OR ROM64_INSTR_PT(571) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(583) OR ROM64_INSTR_PT(584)
     OR ROM64_INSTR_PT(588) OR ROM64_INSTR_PT(592)
     OR ROM64_INSTR_PT(595) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(600) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(609) OR ROM64_INSTR_PT(612)
     OR ROM64_INSTR_PT(613) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(623)
     OR ROM64_INSTR_PT(628) OR ROM64_INSTR_PT(633)
     OR ROM64_INSTR_PT(636) OR ROM64_INSTR_PT(637)
     OR ROM64_INSTR_PT(639) OR ROM64_INSTR_PT(642)
     OR ROM64_INSTR_PT(644) OR ROM64_INSTR_PT(646)
     OR ROM64_INSTR_PT(649) OR ROM64_INSTR_PT(666)
     OR ROM64_INSTR_PT(678) OR ROM64_INSTR_PT(682)
     OR ROM64_INSTR_PT(691) OR ROM64_INSTR_PT(693)
     OR ROM64_INSTR_PT(703) OR ROM64_INSTR_PT(739)
     OR ROM64_INSTR_PT(744) OR ROM64_INSTR_PT(753)
     OR ROM64_INSTR_PT(761) OR ROM64_INSTR_PT(769)
     OR ROM64_INSTR_PT(776) OR ROM64_INSTR_PT(805)
     OR ROM64_INSTR_PT(823) OR ROM64_INSTR_PT(856)
     OR ROM64_INSTR_PT(864) OR ROM64_INSTR_PT(870)
    );
MQQ906:TEMPLATE(15) <= 
    (ROM64_INSTR_PT(9) OR ROM64_INSTR_PT(15)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(53)
     OR ROM64_INSTR_PT(57) OR ROM64_INSTR_PT(71)
     OR ROM64_INSTR_PT(77) OR ROM64_INSTR_PT(80)
     OR ROM64_INSTR_PT(83) OR ROM64_INSTR_PT(89)
     OR ROM64_INSTR_PT(92) OR ROM64_INSTR_PT(96)
     OR ROM64_INSTR_PT(106) OR ROM64_INSTR_PT(110)
     OR ROM64_INSTR_PT(114) OR ROM64_INSTR_PT(116)
     OR ROM64_INSTR_PT(121) OR ROM64_INSTR_PT(122)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(148)
     OR ROM64_INSTR_PT(158) OR ROM64_INSTR_PT(162)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(170)
     OR ROM64_INSTR_PT(173) OR ROM64_INSTR_PT(174)
     OR ROM64_INSTR_PT(175) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(211) OR ROM64_INSTR_PT(213)
     OR ROM64_INSTR_PT(214) OR ROM64_INSTR_PT(218)
     OR ROM64_INSTR_PT(219) OR ROM64_INSTR_PT(222)
     OR ROM64_INSTR_PT(236) OR ROM64_INSTR_PT(240)
     OR ROM64_INSTR_PT(272) OR ROM64_INSTR_PT(273)
     OR ROM64_INSTR_PT(278) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(294) OR ROM64_INSTR_PT(299)
     OR ROM64_INSTR_PT(311) OR ROM64_INSTR_PT(350)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(358)
     OR ROM64_INSTR_PT(363) OR ROM64_INSTR_PT(370)
     OR ROM64_INSTR_PT(371) OR ROM64_INSTR_PT(396)
     OR ROM64_INSTR_PT(399) OR ROM64_INSTR_PT(408)
     OR ROM64_INSTR_PT(416) OR ROM64_INSTR_PT(417)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(425)
     OR ROM64_INSTR_PT(429) OR ROM64_INSTR_PT(433)
     OR ROM64_INSTR_PT(435) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(442) OR ROM64_INSTR_PT(443)
     OR ROM64_INSTR_PT(451) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(461) OR ROM64_INSTR_PT(466)
     OR ROM64_INSTR_PT(474) OR ROM64_INSTR_PT(480)
     OR ROM64_INSTR_PT(506) OR ROM64_INSTR_PT(508)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(532) OR ROM64_INSTR_PT(537)
     OR ROM64_INSTR_PT(562) OR ROM64_INSTR_PT(564)
     OR ROM64_INSTR_PT(581) OR ROM64_INSTR_PT(582)
     OR ROM64_INSTR_PT(585) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(599) OR ROM64_INSTR_PT(603)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(613)
     OR ROM64_INSTR_PT(614) OR ROM64_INSTR_PT(626)
     OR ROM64_INSTR_PT(659) OR ROM64_INSTR_PT(664)
     OR ROM64_INSTR_PT(691) OR ROM64_INSTR_PT(695)
     OR ROM64_INSTR_PT(716) OR ROM64_INSTR_PT(731)
     OR ROM64_INSTR_PT(832) OR ROM64_INSTR_PT(834)
     OR ROM64_INSTR_PT(846) OR ROM64_INSTR_PT(854)
    );
MQQ907:TEMPLATE(16) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(10)
     OR ROM64_INSTR_PT(17) OR ROM64_INSTR_PT(20)
     OR ROM64_INSTR_PT(21) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(49)
     OR ROM64_INSTR_PT(55) OR ROM64_INSTR_PT(64)
     OR ROM64_INSTR_PT(75) OR ROM64_INSTR_PT(77)
     OR ROM64_INSTR_PT(80) OR ROM64_INSTR_PT(83)
     OR ROM64_INSTR_PT(89) OR ROM64_INSTR_PT(96)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(99)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(106)
     OR ROM64_INSTR_PT(110) OR ROM64_INSTR_PT(113)
     OR ROM64_INSTR_PT(114) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(121)
     OR ROM64_INSTR_PT(127) OR ROM64_INSTR_PT(171)
     OR ROM64_INSTR_PT(175) OR ROM64_INSTR_PT(188)
     OR ROM64_INSTR_PT(191) OR ROM64_INSTR_PT(199)
     OR ROM64_INSTR_PT(208) OR ROM64_INSTR_PT(214)
     OR ROM64_INSTR_PT(217) OR ROM64_INSTR_PT(218)
     OR ROM64_INSTR_PT(223) OR ROM64_INSTR_PT(226)
     OR ROM64_INSTR_PT(252) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(257) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(274)
     OR ROM64_INSTR_PT(275) OR ROM64_INSTR_PT(280)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(286)
     OR ROM64_INSTR_PT(315) OR ROM64_INSTR_PT(322)
     OR ROM64_INSTR_PT(331) OR ROM64_INSTR_PT(349)
     OR ROM64_INSTR_PT(363) OR ROM64_INSTR_PT(369)
     OR ROM64_INSTR_PT(371) OR ROM64_INSTR_PT(375)
     OR ROM64_INSTR_PT(391) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(404)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(422)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(437)
     OR ROM64_INSTR_PT(448) OR ROM64_INSTR_PT(466)
     OR ROM64_INSTR_PT(472) OR ROM64_INSTR_PT(481)
     OR ROM64_INSTR_PT(505) OR ROM64_INSTR_PT(521)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(525)
     OR ROM64_INSTR_PT(538) OR ROM64_INSTR_PT(540)
     OR ROM64_INSTR_PT(558) OR ROM64_INSTR_PT(563)
     OR ROM64_INSTR_PT(569) OR ROM64_INSTR_PT(582)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(595)
     OR ROM64_INSTR_PT(596) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(598) OR ROM64_INSTR_PT(600)
     OR ROM64_INSTR_PT(608) OR ROM64_INSTR_PT(613)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(629)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(644)
     OR ROM64_INSTR_PT(744) OR ROM64_INSTR_PT(769)
     OR ROM64_INSTR_PT(776) OR ROM64_INSTR_PT(870)
    );
MQQ908:TEMPLATE(17) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(17)
     OR ROM64_INSTR_PT(20) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(34) OR ROM64_INSTR_PT(38)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(43)
     OR ROM64_INSTR_PT(49) OR ROM64_INSTR_PT(55)
     OR ROM64_INSTR_PT(61) OR ROM64_INSTR_PT(70)
     OR ROM64_INSTR_PT(77) OR ROM64_INSTR_PT(78)
     OR ROM64_INSTR_PT(80) OR ROM64_INSTR_PT(86)
     OR ROM64_INSTR_PT(89) OR ROM64_INSTR_PT(90)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(99)
     OR ROM64_INSTR_PT(102) OR ROM64_INSTR_PT(104)
     OR ROM64_INSTR_PT(106) OR ROM64_INSTR_PT(111)
     OR ROM64_INSTR_PT(114) OR ROM64_INSTR_PT(118)
     OR ROM64_INSTR_PT(121) OR ROM64_INSTR_PT(127)
     OR ROM64_INSTR_PT(144) OR ROM64_INSTR_PT(168)
     OR ROM64_INSTR_PT(173) OR ROM64_INSTR_PT(175)
     OR ROM64_INSTR_PT(186) OR ROM64_INSTR_PT(188)
     OR ROM64_INSTR_PT(191) OR ROM64_INSTR_PT(199)
     OR ROM64_INSTR_PT(208) OR ROM64_INSTR_PT(215)
     OR ROM64_INSTR_PT(219) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(226) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(252) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(257) OR ROM64_INSTR_PT(270)
     OR ROM64_INSTR_PT(271) OR ROM64_INSTR_PT(274)
     OR ROM64_INSTR_PT(277) OR ROM64_INSTR_PT(280)
     OR ROM64_INSTR_PT(282) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(286) OR ROM64_INSTR_PT(287)
     OR ROM64_INSTR_PT(293) OR ROM64_INSTR_PT(302)
     OR ROM64_INSTR_PT(305) OR ROM64_INSTR_PT(322)
     OR ROM64_INSTR_PT(329) OR ROM64_INSTR_PT(331)
     OR ROM64_INSTR_PT(343) OR ROM64_INSTR_PT(349)
     OR ROM64_INSTR_PT(361) OR ROM64_INSTR_PT(364)
     OR ROM64_INSTR_PT(369) OR ROM64_INSTR_PT(383)
     OR ROM64_INSTR_PT(385) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(406)
     OR ROM64_INSTR_PT(408) OR ROM64_INSTR_PT(410)
     OR ROM64_INSTR_PT(420) OR ROM64_INSTR_PT(422)
     OR ROM64_INSTR_PT(424) OR ROM64_INSTR_PT(427)
     OR ROM64_INSTR_PT(448) OR ROM64_INSTR_PT(466)
     OR ROM64_INSTR_PT(472) OR ROM64_INSTR_PT(478)
     OR ROM64_INSTR_PT(480) OR ROM64_INSTR_PT(481)
     OR ROM64_INSTR_PT(482) OR ROM64_INSTR_PT(483)
     OR ROM64_INSTR_PT(484) OR ROM64_INSTR_PT(485)
     OR ROM64_INSTR_PT(493) OR ROM64_INSTR_PT(495)
     OR ROM64_INSTR_PT(498) OR ROM64_INSTR_PT(508)
     OR ROM64_INSTR_PT(511) OR ROM64_INSTR_PT(522)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(534)
     OR ROM64_INSTR_PT(535) OR ROM64_INSTR_PT(536)
     OR ROM64_INSTR_PT(538) OR ROM64_INSTR_PT(548)
     OR ROM64_INSTR_PT(549) OR ROM64_INSTR_PT(552)
     OR ROM64_INSTR_PT(555) OR ROM64_INSTR_PT(563)
     OR ROM64_INSTR_PT(575) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(583) OR ROM64_INSTR_PT(584)
     OR ROM64_INSTR_PT(588) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(599)
     OR ROM64_INSTR_PT(603) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(612) OR ROM64_INSTR_PT(613)
     OR ROM64_INSTR_PT(614) OR ROM64_INSTR_PT(633)
     OR ROM64_INSTR_PT(637) OR ROM64_INSTR_PT(639)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(644)
     OR ROM64_INSTR_PT(646) OR ROM64_INSTR_PT(666)
     OR ROM64_INSTR_PT(678) OR ROM64_INSTR_PT(682)
     OR ROM64_INSTR_PT(703) OR ROM64_INSTR_PT(870)
    );
MQQ909:TEMPLATE(18) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(20)
     OR ROM64_INSTR_PT(21) OR ROM64_INSTR_PT(39)
     OR ROM64_INSTR_PT(49) OR ROM64_INSTR_PT(77)
     OR ROM64_INSTR_PT(80) OR ROM64_INSTR_PT(89)
     OR ROM64_INSTR_PT(97) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(106) OR ROM64_INSTR_PT(110)
     OR ROM64_INSTR_PT(114) OR ROM64_INSTR_PT(118)
     OR ROM64_INSTR_PT(172) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(273)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(397) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(427)
     OR ROM64_INSTR_PT(466) OR ROM64_INSTR_PT(472)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(538)
     OR ROM64_INSTR_PT(544) OR ROM64_INSTR_PT(563)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(733)
    );
MQQ910:TEMPLATE(19) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(15)
     OR ROM64_INSTR_PT(18) OR ROM64_INSTR_PT(20)
     OR ROM64_INSTR_PT(21) OR ROM64_INSTR_PT(25)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(42)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(49)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(57)
     OR ROM64_INSTR_PT(73) OR ROM64_INSTR_PT(77)
     OR ROM64_INSTR_PT(80) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(97) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(106)
     OR ROM64_INSTR_PT(109) OR ROM64_INSTR_PT(118)
     OR ROM64_INSTR_PT(128) OR ROM64_INSTR_PT(145)
     OR ROM64_INSTR_PT(157) OR ROM64_INSTR_PT(168)
     OR ROM64_INSTR_PT(182) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(205) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(219)
     OR ROM64_INSTR_PT(223) OR ROM64_INSTR_PT(236)
     OR ROM64_INSTR_PT(244) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(254) OR ROM64_INSTR_PT(262)
     OR ROM64_INSTR_PT(269) OR ROM64_INSTR_PT(272)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(280)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(290) OR ROM64_INSTR_PT(308)
     OR ROM64_INSTR_PT(325) OR ROM64_INSTR_PT(348)
     OR ROM64_INSTR_PT(361) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(387) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(397) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(406) OR ROM64_INSTR_PT(409)
     OR ROM64_INSTR_PT(419) OR ROM64_INSTR_PT(422)
     OR ROM64_INSTR_PT(425) OR ROM64_INSTR_PT(427)
     OR ROM64_INSTR_PT(429) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(439) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(451) OR ROM64_INSTR_PT(454)
     OR ROM64_INSTR_PT(455) OR ROM64_INSTR_PT(460)
     OR ROM64_INSTR_PT(466) OR ROM64_INSTR_PT(472)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(510) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(532) OR ROM64_INSTR_PT(538)
     OR ROM64_INSTR_PT(539) OR ROM64_INSTR_PT(542)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(570) OR ROM64_INSTR_PT(577)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(582)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(611) OR ROM64_INSTR_PT(616)
     OR ROM64_INSTR_PT(619) OR ROM64_INSTR_PT(636)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(643)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(733)
     OR ROM64_INSTR_PT(736) OR ROM64_INSTR_PT(770)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(823)
     OR ROM64_INSTR_PT(824));
MQQ911:TEMPLATE(20) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(13)
     OR ROM64_INSTR_PT(18) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(35) OR ROM64_INSTR_PT(36)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(42)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(49)
     OR ROM64_INSTR_PT(56) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(162) OR ROM64_INSTR_PT(196)
     OR ROM64_INSTR_PT(216) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(236) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(262)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(280)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(308) OR ROM64_INSTR_PT(325)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(365)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(425)
     OR ROM64_INSTR_PT(426) OR ROM64_INSTR_PT(427)
     OR ROM64_INSTR_PT(429) OR ROM64_INSTR_PT(435)
     OR ROM64_INSTR_PT(439) OR ROM64_INSTR_PT(451)
     OR ROM64_INSTR_PT(454) OR ROM64_INSTR_PT(455)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(466) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(488) OR ROM64_INSTR_PT(507)
     OR ROM64_INSTR_PT(517) OR ROM64_INSTR_PT(520)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(538)
     OR ROM64_INSTR_PT(542) OR ROM64_INSTR_PT(544)
     OR ROM64_INSTR_PT(564) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(586)
     OR ROM64_INSTR_PT(587) OR ROM64_INSTR_PT(589)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(619) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(681)
     OR ROM64_INSTR_PT(693) OR ROM64_INSTR_PT(721)
     OR ROM64_INSTR_PT(728) OR ROM64_INSTR_PT(735)
     OR ROM64_INSTR_PT(738) OR ROM64_INSTR_PT(770)
     OR ROM64_INSTR_PT(811) OR ROM64_INSTR_PT(823)
    );
MQQ912:TEMPLATE(21) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(6)
     OR ROM64_INSTR_PT(9) OR ROM64_INSTR_PT(10)
     OR ROM64_INSTR_PT(11) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(25)
     OR ROM64_INSTR_PT(36) OR ROM64_INSTR_PT(39)
     OR ROM64_INSTR_PT(43) OR ROM64_INSTR_PT(58)
     OR ROM64_INSTR_PT(70) OR ROM64_INSTR_PT(71)
     OR ROM64_INSTR_PT(76) OR ROM64_INSTR_PT(78)
     OR ROM64_INSTR_PT(83) OR ROM64_INSTR_PT(86)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(96)
     OR ROM64_INSTR_PT(97) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(117) OR ROM64_INSTR_PT(118)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(148)
     OR ROM64_INSTR_PT(154) OR ROM64_INSTR_PT(168)
     OR ROM64_INSTR_PT(172) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(182) OR ROM64_INSTR_PT(184)
     OR ROM64_INSTR_PT(188) OR ROM64_INSTR_PT(194)
     OR ROM64_INSTR_PT(201) OR ROM64_INSTR_PT(202)
     OR ROM64_INSTR_PT(205) OR ROM64_INSTR_PT(214)
     OR ROM64_INSTR_PT(216) OR ROM64_INSTR_PT(219)
     OR ROM64_INSTR_PT(222) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(245) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(257) OR ROM64_INSTR_PT(258)
     OR ROM64_INSTR_PT(260) OR ROM64_INSTR_PT(261)
     OR ROM64_INSTR_PT(264) OR ROM64_INSTR_PT(268)
     OR ROM64_INSTR_PT(271) OR ROM64_INSTR_PT(273)
     OR ROM64_INSTR_PT(275) OR ROM64_INSTR_PT(277)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(298) OR ROM64_INSTR_PT(299)
     OR ROM64_INSTR_PT(312) OR ROM64_INSTR_PT(315)
     OR ROM64_INSTR_PT(348) OR ROM64_INSTR_PT(361)
     OR ROM64_INSTR_PT(363) OR ROM64_INSTR_PT(365)
     OR ROM64_INSTR_PT(371) OR ROM64_INSTR_PT(375)
     OR ROM64_INSTR_PT(387) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(391) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(404)
     OR ROM64_INSTR_PT(406) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(424)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(434) OR ROM64_INSTR_PT(437)
     OR ROM64_INSTR_PT(438) OR ROM64_INSTR_PT(457)
     OR ROM64_INSTR_PT(458) OR ROM64_INSTR_PT(463)
     OR ROM64_INSTR_PT(497) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(505) OR ROM64_INSTR_PT(509)
     OR ROM64_INSTR_PT(510) OR ROM64_INSTR_PT(511)
     OR ROM64_INSTR_PT(520) OR ROM64_INSTR_PT(521)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(525)
     OR ROM64_INSTR_PT(530) OR ROM64_INSTR_PT(531)
     OR ROM64_INSTR_PT(535) OR ROM64_INSTR_PT(538)
     OR ROM64_INSTR_PT(540) OR ROM64_INSTR_PT(544)
     OR ROM64_INSTR_PT(545) OR ROM64_INSTR_PT(549)
     OR ROM64_INSTR_PT(558) OR ROM64_INSTR_PT(569)
     OR ROM64_INSTR_PT(570) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(584)
     OR ROM64_INSTR_PT(588) OR ROM64_INSTR_PT(592)
     OR ROM64_INSTR_PT(595) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(598) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(623)
     OR ROM64_INSTR_PT(628) OR ROM64_INSTR_PT(629)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(728)
     OR ROM64_INSTR_PT(735) OR ROM64_INSTR_PT(738)
     OR ROM64_INSTR_PT(822));
MQQ913:TEMPLATE(22) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(8)
     OR ROM64_INSTR_PT(9) OR ROM64_INSTR_PT(11)
     OR ROM64_INSTR_PT(13) OR ROM64_INSTR_PT(15)
     OR ROM64_INSTR_PT(18) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(25)
     OR ROM64_INSTR_PT(30) OR ROM64_INSTR_PT(36)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(43)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(56)
     OR ROM64_INSTR_PT(57) OR ROM64_INSTR_PT(71)
     OR ROM64_INSTR_PT(73) OR ROM64_INSTR_PT(76)
     OR ROM64_INSTR_PT(78) OR ROM64_INSTR_PT(93)
     OR ROM64_INSTR_PT(97) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(113)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(121)
     OR ROM64_INSTR_PT(128) OR ROM64_INSTR_PT(133)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(148)
     OR ROM64_INSTR_PT(155) OR ROM64_INSTR_PT(157)
     OR ROM64_INSTR_PT(162) OR ROM64_INSTR_PT(164)
     OR ROM64_INSTR_PT(171) OR ROM64_INSTR_PT(172)
     OR ROM64_INSTR_PT(175) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(184) OR ROM64_INSTR_PT(188)
     OR ROM64_INSTR_PT(196) OR ROM64_INSTR_PT(201)
     OR ROM64_INSTR_PT(202) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(206) OR ROM64_INSTR_PT(211)
     OR ROM64_INSTR_PT(216) OR ROM64_INSTR_PT(218)
     OR ROM64_INSTR_PT(222) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(244) OR ROM64_INSTR_PT(245)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(257)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(272)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(280)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(298)
     OR ROM64_INSTR_PT(299) OR ROM64_INSTR_PT(312)
     OR ROM64_INSTR_PT(325) OR ROM64_INSTR_PT(353)
     OR ROM64_INSTR_PT(365) OR ROM64_INSTR_PT(372)
     OR ROM64_INSTR_PT(381) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(414) OR ROM64_INSTR_PT(426)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(434)
     OR ROM64_INSTR_PT(438) OR ROM64_INSTR_PT(439)
     OR ROM64_INSTR_PT(440) OR ROM64_INSTR_PT(443)
     OR ROM64_INSTR_PT(454) OR ROM64_INSTR_PT(455)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(457)
     OR ROM64_INSTR_PT(458) OR ROM64_INSTR_PT(460)
     OR ROM64_INSTR_PT(463) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(481) OR ROM64_INSTR_PT(488)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(497)
     OR ROM64_INSTR_PT(503) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(514)
     OR ROM64_INSTR_PT(519) OR ROM64_INSTR_PT(520)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(532)
     OR ROM64_INSTR_PT(538) OR ROM64_INSTR_PT(539)
     OR ROM64_INSTR_PT(540) OR ROM64_INSTR_PT(544)
     OR ROM64_INSTR_PT(545) OR ROM64_INSTR_PT(553)
     OR ROM64_INSTR_PT(554) OR ROM64_INSTR_PT(566)
     OR ROM64_INSTR_PT(568) OR ROM64_INSTR_PT(576)
     OR ROM64_INSTR_PT(581) OR ROM64_INSTR_PT(582)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(586)
     OR ROM64_INSTR_PT(587) OR ROM64_INSTR_PT(589)
     OR ROM64_INSTR_PT(592) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(598)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(607)
     OR ROM64_INSTR_PT(611) OR ROM64_INSTR_PT(613)
     OR ROM64_INSTR_PT(617) OR ROM64_INSTR_PT(625)
     OR ROM64_INSTR_PT(628) OR ROM64_INSTR_PT(636)
     OR ROM64_INSTR_PT(643) OR ROM64_INSTR_PT(655)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(681)
     OR ROM64_INSTR_PT(698) OR ROM64_INSTR_PT(713)
     OR ROM64_INSTR_PT(723) OR ROM64_INSTR_PT(724)
     OR ROM64_INSTR_PT(728) OR ROM64_INSTR_PT(733)
     OR ROM64_INSTR_PT(735) OR ROM64_INSTR_PT(738)
     OR ROM64_INSTR_PT(822) OR ROM64_INSTR_PT(824)
     OR ROM64_INSTR_PT(846) OR ROM64_INSTR_PT(854)
    );
MQQ914:TEMPLATE(23) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(6)
     OR ROM64_INSTR_PT(13) OR ROM64_INSTR_PT(25)
     OR ROM64_INSTR_PT(36) OR ROM64_INSTR_PT(39)
     OR ROM64_INSTR_PT(56) OR ROM64_INSTR_PT(57)
     OR ROM64_INSTR_PT(73) OR ROM64_INSTR_PT(89)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(100) OR ROM64_INSTR_PT(101)
     OR ROM64_INSTR_PT(110) OR ROM64_INSTR_PT(114)
     OR ROM64_INSTR_PT(124) OR ROM64_INSTR_PT(128)
     OR ROM64_INSTR_PT(137) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(157) OR ROM64_INSTR_PT(162)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(184) OR ROM64_INSTR_PT(194)
     OR ROM64_INSTR_PT(201) OR ROM64_INSTR_PT(202)
     OR ROM64_INSTR_PT(203) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(216) OR ROM64_INSTR_PT(218)
     OR ROM64_INSTR_PT(219) OR ROM64_INSTR_PT(229)
     OR ROM64_INSTR_PT(230) OR ROM64_INSTR_PT(244)
     OR ROM64_INSTR_PT(245) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(263)
     OR ROM64_INSTR_PT(277) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(285) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(312) OR ROM64_INSTR_PT(319)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(361)
     OR ROM64_INSTR_PT(365) OR ROM64_INSTR_PT(372)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(388) OR ROM64_INSTR_PT(395)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(406) OR ROM64_INSTR_PT(413)
     OR ROM64_INSTR_PT(426) OR ROM64_INSTR_PT(434)
     OR ROM64_INSTR_PT(438) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(457)
     OR ROM64_INSTR_PT(458) OR ROM64_INSTR_PT(460)
     OR ROM64_INSTR_PT(467) OR ROM64_INSTR_PT(473)
     OR ROM64_INSTR_PT(475) OR ROM64_INSTR_PT(488)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(517) OR ROM64_INSTR_PT(520)
     OR ROM64_INSTR_PT(531) OR ROM64_INSTR_PT(535)
     OR ROM64_INSTR_PT(538) OR ROM64_INSTR_PT(539)
     OR ROM64_INSTR_PT(545) OR ROM64_INSTR_PT(546)
     OR ROM64_INSTR_PT(549) OR ROM64_INSTR_PT(553)
     OR ROM64_INSTR_PT(554) OR ROM64_INSTR_PT(559)
     OR ROM64_INSTR_PT(563) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(575) OR ROM64_INSTR_PT(582)
     OR ROM64_INSTR_PT(592) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(611)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(623) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(636) OR ROM64_INSTR_PT(643)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(693)
     OR ROM64_INSTR_PT(717) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(728)
     OR ROM64_INSTR_PT(733) OR ROM64_INSTR_PT(735)
     OR ROM64_INSTR_PT(738) OR ROM64_INSTR_PT(822)
     OR ROM64_INSTR_PT(824) OR ROM64_INSTR_PT(846)
    );
MQQ915:TEMPLATE(24) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(11)
     OR ROM64_INSTR_PT(14) OR ROM64_INSTR_PT(30)
     OR ROM64_INSTR_PT(36) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(51)
     OR ROM64_INSTR_PT(77) OR ROM64_INSTR_PT(80)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(100) OR ROM64_INSTR_PT(105)
     OR ROM64_INSTR_PT(106) OR ROM64_INSTR_PT(115)
     OR ROM64_INSTR_PT(124) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(143)
     OR ROM64_INSTR_PT(153) OR ROM64_INSTR_PT(158)
     OR ROM64_INSTR_PT(170) OR ROM64_INSTR_PT(172)
     OR ROM64_INSTR_PT(184) OR ROM64_INSTR_PT(185)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(202)
     OR ROM64_INSTR_PT(204) OR ROM64_INSTR_PT(216)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(229)
     OR ROM64_INSTR_PT(230) OR ROM64_INSTR_PT(241)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(258)
     OR ROM64_INSTR_PT(260) OR ROM64_INSTR_PT(261)
     OR ROM64_INSTR_PT(262) OR ROM64_INSTR_PT(263)
     OR ROM64_INSTR_PT(277) OR ROM64_INSTR_PT(278)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(285)
     OR ROM64_INSTR_PT(294) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(308) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(319) OR ROM64_INSTR_PT(348)
     OR ROM64_INSTR_PT(365) OR ROM64_INSTR_PT(366)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(387)
     OR ROM64_INSTR_PT(394) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(428) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(432) OR ROM64_INSTR_PT(433)
     OR ROM64_INSTR_PT(434) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(453) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(496) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(512)
     OR ROM64_INSTR_PT(520) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(531) OR ROM64_INSTR_PT(535)
     OR ROM64_INSTR_PT(544) OR ROM64_INSTR_PT(545)
     OR ROM64_INSTR_PT(546) OR ROM64_INSTR_PT(549)
     OR ROM64_INSTR_PT(557) OR ROM64_INSTR_PT(559)
     OR ROM64_INSTR_PT(564) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(580)
     OR ROM64_INSTR_PT(582) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(606)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(619) OR ROM64_INSTR_PT(623)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(645) OR ROM64_INSTR_PT(663)
     OR ROM64_INSTR_PT(693) OR ROM64_INSTR_PT(705)
     OR ROM64_INSTR_PT(736) OR ROM64_INSTR_PT(753)
     OR ROM64_INSTR_PT(770) OR ROM64_INSTR_PT(822)
     OR ROM64_INSTR_PT(846));
MQQ916:TEMPLATE(25) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(6)
     OR ROM64_INSTR_PT(13) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(25) OR ROM64_INSTR_PT(36)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(56)
     OR ROM64_INSTR_PT(57) OR ROM64_INSTR_PT(73)
     OR ROM64_INSTR_PT(97) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(118)
     OR ROM64_INSTR_PT(125) OR ROM64_INSTR_PT(128)
     OR ROM64_INSTR_PT(134) OR ROM64_INSTR_PT(143)
     OR ROM64_INSTR_PT(155) OR ROM64_INSTR_PT(157)
     OR ROM64_INSTR_PT(158) OR ROM64_INSTR_PT(162)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(170)
     OR ROM64_INSTR_PT(172) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(182) OR ROM64_INSTR_PT(184)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(196)
     OR ROM64_INSTR_PT(202) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(206) OR ROM64_INSTR_PT(216)
     OR ROM64_INSTR_PT(219) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(244) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(260) OR ROM64_INSTR_PT(261)
     OR ROM64_INSTR_PT(277) OR ROM64_INSTR_PT(278)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(294) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(339) OR ROM64_INSTR_PT(348)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(361)
     OR ROM64_INSTR_PT(365) OR ROM64_INSTR_PT(366)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(387) OR ROM64_INSTR_PT(395)
     OR ROM64_INSTR_PT(397) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(405) OR ROM64_INSTR_PT(406)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(426)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(433) OR ROM64_INSTR_PT(434)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(460) OR ROM64_INSTR_PT(466)
     OR ROM64_INSTR_PT(467) OR ROM64_INSTR_PT(473)
     OR ROM64_INSTR_PT(475) OR ROM64_INSTR_PT(488)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(506) OR ROM64_INSTR_PT(507)
     OR ROM64_INSTR_PT(517) OR ROM64_INSTR_PT(520)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(531) OR ROM64_INSTR_PT(535)
     OR ROM64_INSTR_PT(539) OR ROM64_INSTR_PT(542)
     OR ROM64_INSTR_PT(545) OR ROM64_INSTR_PT(549)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(557) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(575) OR ROM64_INSTR_PT(576)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(584)
     OR ROM64_INSTR_PT(585) OR ROM64_INSTR_PT(592)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(611)
     OR ROM64_INSTR_PT(617) OR ROM64_INSTR_PT(626)
     OR ROM64_INSTR_PT(632) OR ROM64_INSTR_PT(636)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(643)
     OR ROM64_INSTR_PT(649) OR ROM64_INSTR_PT(655)
     OR ROM64_INSTR_PT(664) OR ROM64_INSTR_PT(693)
     OR ROM64_INSTR_PT(702) OR ROM64_INSTR_PT(713)
     OR ROM64_INSTR_PT(736) OR ROM64_INSTR_PT(739)
     OR ROM64_INSTR_PT(753) OR ROM64_INSTR_PT(798)
     OR ROM64_INSTR_PT(822) OR ROM64_INSTR_PT(823)
     OR ROM64_INSTR_PT(824) OR ROM64_INSTR_PT(832)
    );
MQQ917:TEMPLATE(26) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(7)
     OR ROM64_INSTR_PT(9) OR ROM64_INSTR_PT(11)
     OR ROM64_INSTR_PT(14) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(25)
     OR ROM64_INSTR_PT(30) OR ROM64_INSTR_PT(35)
     OR ROM64_INSTR_PT(36) OR ROM64_INSTR_PT(38)
     OR ROM64_INSTR_PT(41) OR ROM64_INSTR_PT(43)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(50)
     OR ROM64_INSTR_PT(51) OR ROM64_INSTR_PT(52)
     OR ROM64_INSTR_PT(56) OR ROM64_INSTR_PT(57)
     OR ROM64_INSTR_PT(58) OR ROM64_INSTR_PT(61)
     OR ROM64_INSTR_PT(68) OR ROM64_INSTR_PT(69)
     OR ROM64_INSTR_PT(70) OR ROM64_INSTR_PT(71)
     OR ROM64_INSTR_PT(73) OR ROM64_INSTR_PT(76)
     OR ROM64_INSTR_PT(78) OR ROM64_INSTR_PT(82)
     OR ROM64_INSTR_PT(83) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(86) OR ROM64_INSTR_PT(90)
     OR ROM64_INSTR_PT(92) OR ROM64_INSTR_PT(93)
     OR ROM64_INSTR_PT(95) OR ROM64_INSTR_PT(97)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(100)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(102)
     OR ROM64_INSTR_PT(105) OR ROM64_INSTR_PT(108)
     OR ROM64_INSTR_PT(109) OR ROM64_INSTR_PT(115)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(124)
     OR ROM64_INSTR_PT(128) OR ROM64_INSTR_PT(132)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(143)
     OR ROM64_INSTR_PT(144) OR ROM64_INSTR_PT(145)
     OR ROM64_INSTR_PT(148) OR ROM64_INSTR_PT(153)
     OR ROM64_INSTR_PT(154) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(157) OR ROM64_INSTR_PT(158)
     OR ROM64_INSTR_PT(162) OR ROM64_INSTR_PT(169)
     OR ROM64_INSTR_PT(172) OR ROM64_INSTR_PT(174)
     OR ROM64_INSTR_PT(177) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(181) OR ROM64_INSTR_PT(183)
     OR ROM64_INSTR_PT(185) OR ROM64_INSTR_PT(186)
     OR ROM64_INSTR_PT(188) OR ROM64_INSTR_PT(194)
     OR ROM64_INSTR_PT(196) OR ROM64_INSTR_PT(201)
     OR ROM64_INSTR_PT(203) OR ROM64_INSTR_PT(204)
     OR ROM64_INSTR_PT(205) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(215) OR ROM64_INSTR_PT(216)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(222)
     OR ROM64_INSTR_PT(223) OR ROM64_INSTR_PT(226)
     OR ROM64_INSTR_PT(233) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(241) OR ROM64_INSTR_PT(243)
     OR ROM64_INSTR_PT(244) OR ROM64_INSTR_PT(245)
     OR ROM64_INSTR_PT(249) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(254) OR ROM64_INSTR_PT(257)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(263)
     OR ROM64_INSTR_PT(264) OR ROM64_INSTR_PT(265)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(269)
     OR ROM64_INSTR_PT(270) OR ROM64_INSTR_PT(271)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(275)
     OR ROM64_INSTR_PT(276) OR ROM64_INSTR_PT(277)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(282)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(285) OR ROM64_INSTR_PT(287)
     OR ROM64_INSTR_PT(290) OR ROM64_INSTR_PT(293)
     OR ROM64_INSTR_PT(294) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(298) OR ROM64_INSTR_PT(299)
     OR ROM64_INSTR_PT(302) OR ROM64_INSTR_PT(305)
     OR ROM64_INSTR_PT(308) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(312) OR ROM64_INSTR_PT(315)
     OR ROM64_INSTR_PT(319) OR ROM64_INSTR_PT(339)
     OR ROM64_INSTR_PT(348) OR ROM64_INSTR_PT(350)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(355)
     OR ROM64_INSTR_PT(358) OR ROM64_INSTR_PT(364)
     OR ROM64_INSTR_PT(365) OR ROM64_INSTR_PT(367)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(374)
     OR ROM64_INSTR_PT(375) OR ROM64_INSTR_PT(378)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(383) OR ROM64_INSTR_PT(384)
     OR ROM64_INSTR_PT(385) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(391) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(403)
     OR ROM64_INSTR_PT(404) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(409) OR ROM64_INSTR_PT(410)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(419) OR ROM64_INSTR_PT(424)
     OR ROM64_INSTR_PT(425) OR ROM64_INSTR_PT(426)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(428)
     OR ROM64_INSTR_PT(429) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(432) OR ROM64_INSTR_PT(435)
     OR ROM64_INSTR_PT(437) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(451)
     OR ROM64_INSTR_PT(453) OR ROM64_INSTR_PT(456)
     OR ROM64_INSTR_PT(457) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(460) OR ROM64_INSTR_PT(461)
     OR ROM64_INSTR_PT(463) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(478) OR ROM64_INSTR_PT(481)
     OR ROM64_INSTR_PT(482) OR ROM64_INSTR_PT(484)
     OR ROM64_INSTR_PT(485) OR ROM64_INSTR_PT(488)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(493)
     OR ROM64_INSTR_PT(495) OR ROM64_INSTR_PT(496)
     OR ROM64_INSTR_PT(497) OR ROM64_INSTR_PT(504)
     OR ROM64_INSTR_PT(505) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(510)
     OR ROM64_INSTR_PT(511) OR ROM64_INSTR_PT(512)
     OR ROM64_INSTR_PT(517) OR ROM64_INSTR_PT(520)
     OR ROM64_INSTR_PT(521) OR ROM64_INSTR_PT(522)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(525)
     OR ROM64_INSTR_PT(530) OR ROM64_INSTR_PT(531)
     OR ROM64_INSTR_PT(534) OR ROM64_INSTR_PT(535)
     OR ROM64_INSTR_PT(539) OR ROM64_INSTR_PT(540)
     OR ROM64_INSTR_PT(544) OR ROM64_INSTR_PT(546)
     OR ROM64_INSTR_PT(549) OR ROM64_INSTR_PT(552)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(555) OR ROM64_INSTR_PT(557)
     OR ROM64_INSTR_PT(558) OR ROM64_INSTR_PT(559)
     OR ROM64_INSTR_PT(563) OR ROM64_INSTR_PT(564)
     OR ROM64_INSTR_PT(568) OR ROM64_INSTR_PT(569)
     OR ROM64_INSTR_PT(570) OR ROM64_INSTR_PT(571)
     OR ROM64_INSTR_PT(575) OR ROM64_INSTR_PT(576)
     OR ROM64_INSTR_PT(577) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(582)
     OR ROM64_INSTR_PT(583) OR ROM64_INSTR_PT(584)
     OR ROM64_INSTR_PT(588) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(592) OR ROM64_INSTR_PT(595)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(598)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(609) OR ROM64_INSTR_PT(611)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(616)
     OR ROM64_INSTR_PT(617) OR ROM64_INSTR_PT(618)
     OR ROM64_INSTR_PT(619) OR ROM64_INSTR_PT(623)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(629) OR ROM64_INSTR_PT(632)
     OR ROM64_INSTR_PT(633) OR ROM64_INSTR_PT(636)
     OR ROM64_INSTR_PT(639) OR ROM64_INSTR_PT(642)
     OR ROM64_INSTR_PT(643) OR ROM64_INSTR_PT(655)
     OR ROM64_INSTR_PT(660) OR ROM64_INSTR_PT(663)
     OR ROM64_INSTR_PT(664) OR ROM64_INSTR_PT(666)
     OR ROM64_INSTR_PT(678) OR ROM64_INSTR_PT(695)
     OR ROM64_INSTR_PT(702) OR ROM64_INSTR_PT(713)
     OR ROM64_INSTR_PT(716) OR ROM64_INSTR_PT(717)
     OR ROM64_INSTR_PT(721) OR ROM64_INSTR_PT(722)
     OR ROM64_INSTR_PT(723) OR ROM64_INSTR_PT(724)
     OR ROM64_INSTR_PT(733) OR ROM64_INSTR_PT(736)
     OR ROM64_INSTR_PT(761) OR ROM64_INSTR_PT(770)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(811)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(822)
     OR ROM64_INSTR_PT(824) OR ROM64_INSTR_PT(832)
     OR ROM64_INSTR_PT(834) OR ROM64_INSTR_PT(846)
     OR ROM64_INSTR_PT(855) OR ROM64_INSTR_PT(856)
     OR ROM64_INSTR_PT(858) OR ROM64_INSTR_PT(864)
     OR ROM64_INSTR_PT(870) OR ROM64_INSTR_PT(873)
    );
MQQ918:TEMPLATE(27) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(6)
     OR ROM64_INSTR_PT(7) OR ROM64_INSTR_PT(8)
     OR ROM64_INSTR_PT(9) OR ROM64_INSTR_PT(11)
     OR ROM64_INSTR_PT(15) OR ROM64_INSTR_PT(18)
     OR ROM64_INSTR_PT(21) OR ROM64_INSTR_PT(22)
     OR ROM64_INSTR_PT(35) OR ROM64_INSTR_PT(38)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(45)
     OR ROM64_INSTR_PT(49) OR ROM64_INSTR_PT(52)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(56)
     OR ROM64_INSTR_PT(57) OR ROM64_INSTR_PT(61)
     OR ROM64_INSTR_PT(68) OR ROM64_INSTR_PT(69)
     OR ROM64_INSTR_PT(71) OR ROM64_INSTR_PT(73)
     OR ROM64_INSTR_PT(82) OR ROM64_INSTR_PT(83)
     OR ROM64_INSTR_PT(84) OR ROM64_INSTR_PT(90)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(95)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(101)
     OR ROM64_INSTR_PT(102) OR ROM64_INSTR_PT(108)
     OR ROM64_INSTR_PT(109) OR ROM64_INSTR_PT(113)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(128)
     OR ROM64_INSTR_PT(132) OR ROM64_INSTR_PT(133)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(143)
     OR ROM64_INSTR_PT(144) OR ROM64_INSTR_PT(145)
     OR ROM64_INSTR_PT(148) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(157) OR ROM64_INSTR_PT(158)
     OR ROM64_INSTR_PT(162) OR ROM64_INSTR_PT(164)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(169)
     OR ROM64_INSTR_PT(170) OR ROM64_INSTR_PT(171)
     OR ROM64_INSTR_PT(177) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(181) OR ROM64_INSTR_PT(182)
     OR ROM64_INSTR_PT(183) OR ROM64_INSTR_PT(186)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(196)
     OR ROM64_INSTR_PT(201) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(205) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(211) OR ROM64_INSTR_PT(215)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(219)
     OR ROM64_INSTR_PT(222) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(226) OR ROM64_INSTR_PT(233)
     OR ROM64_INSTR_PT(238) OR ROM64_INSTR_PT(240)
     OR ROM64_INSTR_PT(243) OR ROM64_INSTR_PT(244)
     OR ROM64_INSTR_PT(245) OR ROM64_INSTR_PT(249)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(254)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(264) OR ROM64_INSTR_PT(265)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(269)
     OR ROM64_INSTR_PT(270) OR ROM64_INSTR_PT(272)
     OR ROM64_INSTR_PT(276) OR ROM64_INSTR_PT(278)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(282)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(287) OR ROM64_INSTR_PT(290)
     OR ROM64_INSTR_PT(293) OR ROM64_INSTR_PT(294)
     OR ROM64_INSTR_PT(298) OR ROM64_INSTR_PT(299)
     OR ROM64_INSTR_PT(302) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(312) OR ROM64_INSTR_PT(325)
     OR ROM64_INSTR_PT(339) OR ROM64_INSTR_PT(348)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(361)
     OR ROM64_INSTR_PT(364) OR ROM64_INSTR_PT(366)
     OR ROM64_INSTR_PT(367) OR ROM64_INSTR_PT(372)
     OR ROM64_INSTR_PT(374) OR ROM64_INSTR_PT(375)
     OR ROM64_INSTR_PT(378) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(383) OR ROM64_INSTR_PT(384)
     OR ROM64_INSTR_PT(385) OR ROM64_INSTR_PT(391)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(396)
     OR ROM64_INSTR_PT(397) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(403) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(406) OR ROM64_INSTR_PT(409)
     OR ROM64_INSTR_PT(410) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(419) OR ROM64_INSTR_PT(425)
     OR ROM64_INSTR_PT(426) OR ROM64_INSTR_PT(427)
     OR ROM64_INSTR_PT(428) OR ROM64_INSTR_PT(429)
     OR ROM64_INSTR_PT(430) OR ROM64_INSTR_PT(433)
     OR ROM64_INSTR_PT(435) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(439) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(443) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(451) OR ROM64_INSTR_PT(454)
     OR ROM64_INSTR_PT(455) OR ROM64_INSTR_PT(456)
     OR ROM64_INSTR_PT(457) OR ROM64_INSTR_PT(460)
     OR ROM64_INSTR_PT(467) OR ROM64_INSTR_PT(473)
     OR ROM64_INSTR_PT(475) OR ROM64_INSTR_PT(478)
     OR ROM64_INSTR_PT(481) OR ROM64_INSTR_PT(482)
     OR ROM64_INSTR_PT(484) OR ROM64_INSTR_PT(485)
     OR ROM64_INSTR_PT(488) OR ROM64_INSTR_PT(490)
     OR ROM64_INSTR_PT(495) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(510)
     OR ROM64_INSTR_PT(514) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(522) OR ROM64_INSTR_PT(523)
     OR ROM64_INSTR_PT(525) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(531) OR ROM64_INSTR_PT(532)
     OR ROM64_INSTR_PT(534) OR ROM64_INSTR_PT(539)
     OR ROM64_INSTR_PT(542) OR ROM64_INSTR_PT(552)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(555) OR ROM64_INSTR_PT(557)
     OR ROM64_INSTR_PT(563) OR ROM64_INSTR_PT(564)
     OR ROM64_INSTR_PT(566) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(570) OR ROM64_INSTR_PT(571)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(577)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(581)
     OR ROM64_INSTR_PT(582) OR ROM64_INSTR_PT(583)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(585)
     OR ROM64_INSTR_PT(586) OR ROM64_INSTR_PT(587)
     OR ROM64_INSTR_PT(589) OR ROM64_INSTR_PT(592)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(604)
     OR ROM64_INSTR_PT(607) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(611) OR ROM64_INSTR_PT(616)
     OR ROM64_INSTR_PT(619) OR ROM64_INSTR_PT(625)
     OR ROM64_INSTR_PT(626) OR ROM64_INSTR_PT(629)
     OR ROM64_INSTR_PT(632) OR ROM64_INSTR_PT(633)
     OR ROM64_INSTR_PT(636) OR ROM64_INSTR_PT(639)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(643)
     OR ROM64_INSTR_PT(655) OR ROM64_INSTR_PT(660)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(664)
     OR ROM64_INSTR_PT(666) OR ROM64_INSTR_PT(678)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(698)
     OR ROM64_INSTR_PT(702) OR ROM64_INSTR_PT(713)
     OR ROM64_INSTR_PT(722) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(733)
     OR ROM64_INSTR_PT(736) OR ROM64_INSTR_PT(753)
     OR ROM64_INSTR_PT(761) OR ROM64_INSTR_PT(770)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(811)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(823)
     OR ROM64_INSTR_PT(824) OR ROM64_INSTR_PT(832)
     OR ROM64_INSTR_PT(834) OR ROM64_INSTR_PT(854)
     OR ROM64_INSTR_PT(855) OR ROM64_INSTR_PT(856)
     OR ROM64_INSTR_PT(864) OR ROM64_INSTR_PT(870)
    );
MQQ919:TEMPLATE(28) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(9)
     OR ROM64_INSTR_PT(14) OR ROM64_INSTR_PT(17)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(38) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(51)
     OR ROM64_INSTR_PT(52) OR ROM64_INSTR_PT(56)
     OR ROM64_INSTR_PT(57) OR ROM64_INSTR_PT(61)
     OR ROM64_INSTR_PT(64) OR ROM64_INSTR_PT(68)
     OR ROM64_INSTR_PT(69) OR ROM64_INSTR_PT(70)
     OR ROM64_INSTR_PT(71) OR ROM64_INSTR_PT(73)
     OR ROM64_INSTR_PT(75) OR ROM64_INSTR_PT(82)
     OR ROM64_INSTR_PT(83) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(86) OR ROM64_INSTR_PT(90)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(95)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(99)
     OR ROM64_INSTR_PT(100) OR ROM64_INSTR_PT(101)
     OR ROM64_INSTR_PT(102) OR ROM64_INSTR_PT(105)
     OR ROM64_INSTR_PT(108) OR ROM64_INSTR_PT(113)
     OR ROM64_INSTR_PT(115) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(124) OR ROM64_INSTR_PT(125)
     OR ROM64_INSTR_PT(127) OR ROM64_INSTR_PT(128)
     OR ROM64_INSTR_PT(134) OR ROM64_INSTR_PT(136)
     OR ROM64_INSTR_PT(137) OR ROM64_INSTR_PT(140)
     OR ROM64_INSTR_PT(143) OR ROM64_INSTR_PT(144)
     OR ROM64_INSTR_PT(148) OR ROM64_INSTR_PT(153)
     OR ROM64_INSTR_PT(155) OR ROM64_INSTR_PT(157)
     OR ROM64_INSTR_PT(158) OR ROM64_INSTR_PT(162)
     OR ROM64_INSTR_PT(169) OR ROM64_INSTR_PT(171)
     OR ROM64_INSTR_PT(180) OR ROM64_INSTR_PT(185)
     OR ROM64_INSTR_PT(186) OR ROM64_INSTR_PT(194)
     OR ROM64_INSTR_PT(196) OR ROM64_INSTR_PT(199)
     OR ROM64_INSTR_PT(201) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(204) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(215) OR ROM64_INSTR_PT(217)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(222)
     OR ROM64_INSTR_PT(226) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(241) OR ROM64_INSTR_PT(243)
     OR ROM64_INSTR_PT(244) OR ROM64_INSTR_PT(249)
     OR ROM64_INSTR_PT(252) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(263) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(265) OR ROM64_INSTR_PT(268)
     OR ROM64_INSTR_PT(269) OR ROM64_INSTR_PT(270)
     OR ROM64_INSTR_PT(271) OR ROM64_INSTR_PT(275)
     OR ROM64_INSTR_PT(282) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(284) OR ROM64_INSTR_PT(285)
     OR ROM64_INSTR_PT(287) OR ROM64_INSTR_PT(290)
     OR ROM64_INSTR_PT(293) OR ROM64_INSTR_PT(294)
     OR ROM64_INSTR_PT(297) OR ROM64_INSTR_PT(298)
     OR ROM64_INSTR_PT(299) OR ROM64_INSTR_PT(302)
     OR ROM64_INSTR_PT(305) OR ROM64_INSTR_PT(308)
     OR ROM64_INSTR_PT(311) OR ROM64_INSTR_PT(315)
     OR ROM64_INSTR_PT(319) OR ROM64_INSTR_PT(331)
     OR ROM64_INSTR_PT(339) OR ROM64_INSTR_PT(348)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(364)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(374)
     OR ROM64_INSTR_PT(375) OR ROM64_INSTR_PT(379)
     OR ROM64_INSTR_PT(381) OR ROM64_INSTR_PT(383)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(385)
     OR ROM64_INSTR_PT(391) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(404) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(410) OR ROM64_INSTR_PT(413)
     OR ROM64_INSTR_PT(414) OR ROM64_INSTR_PT(415)
     OR ROM64_INSTR_PT(418) OR ROM64_INSTR_PT(424)
     OR ROM64_INSTR_PT(425) OR ROM64_INSTR_PT(426)
     OR ROM64_INSTR_PT(428) OR ROM64_INSTR_PT(429)
     OR ROM64_INSTR_PT(430) OR ROM64_INSTR_PT(432)
     OR ROM64_INSTR_PT(435) OR ROM64_INSTR_PT(437)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(451) OR ROM64_INSTR_PT(453)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(457)
     OR ROM64_INSTR_PT(460) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(478) OR ROM64_INSTR_PT(481)
     OR ROM64_INSTR_PT(482) OR ROM64_INSTR_PT(484)
     OR ROM64_INSTR_PT(485) OR ROM64_INSTR_PT(488)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(493)
     OR ROM64_INSTR_PT(495) OR ROM64_INSTR_PT(496)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(505)
     OR ROM64_INSTR_PT(506) OR ROM64_INSTR_PT(507)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(511)
     OR ROM64_INSTR_PT(512) OR ROM64_INSTR_PT(517)
     OR ROM64_INSTR_PT(521) OR ROM64_INSTR_PT(522)
     OR ROM64_INSTR_PT(525) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(531) OR ROM64_INSTR_PT(534)
     OR ROM64_INSTR_PT(539) OR ROM64_INSTR_PT(546)
     OR ROM64_INSTR_PT(552) OR ROM64_INSTR_PT(553)
     OR ROM64_INSTR_PT(554) OR ROM64_INSTR_PT(555)
     OR ROM64_INSTR_PT(557) OR ROM64_INSTR_PT(558)
     OR ROM64_INSTR_PT(559) OR ROM64_INSTR_PT(563)
     OR ROM64_INSTR_PT(564) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(569) OR ROM64_INSTR_PT(577)
     OR ROM64_INSTR_PT(579) OR ROM64_INSTR_PT(580)
     OR ROM64_INSTR_PT(582) OR ROM64_INSTR_PT(583)
     OR ROM64_INSTR_PT(588) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(592) OR ROM64_INSTR_PT(595)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(600)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(611) OR ROM64_INSTR_PT(615)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(619)
     OR ROM64_INSTR_PT(623) OR ROM64_INSTR_PT(627)
     OR ROM64_INSTR_PT(629) OR ROM64_INSTR_PT(632)
     OR ROM64_INSTR_PT(633) OR ROM64_INSTR_PT(636)
     OR ROM64_INSTR_PT(639) OR ROM64_INSTR_PT(642)
     OR ROM64_INSTR_PT(643) OR ROM64_INSTR_PT(644)
     OR ROM64_INSTR_PT(655) OR ROM64_INSTR_PT(660)
     OR ROM64_INSTR_PT(664) OR ROM64_INSTR_PT(666)
     OR ROM64_INSTR_PT(678) OR ROM64_INSTR_PT(702)
     OR ROM64_INSTR_PT(713) OR ROM64_INSTR_PT(722)
     OR ROM64_INSTR_PT(728) OR ROM64_INSTR_PT(735)
     OR ROM64_INSTR_PT(736) OR ROM64_INSTR_PT(738)
     OR ROM64_INSTR_PT(739) OR ROM64_INSTR_PT(744)
     OR ROM64_INSTR_PT(761) OR ROM64_INSTR_PT(769)
     OR ROM64_INSTR_PT(770) OR ROM64_INSTR_PT(776)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(811)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(824)
     OR ROM64_INSTR_PT(832) OR ROM64_INSTR_PT(855)
     OR ROM64_INSTR_PT(856) OR ROM64_INSTR_PT(864)
     OR ROM64_INSTR_PT(870));
MQQ920:TEMPLATE(29) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(7)
     OR ROM64_INSTR_PT(8) OR ROM64_INSTR_PT(9)
     OR ROM64_INSTR_PT(11) OR ROM64_INSTR_PT(14)
     OR ROM64_INSTR_PT(15) OR ROM64_INSTR_PT(17)
     OR ROM64_INSTR_PT(18) OR ROM64_INSTR_PT(22)
     OR ROM64_INSTR_PT(25) OR ROM64_INSTR_PT(28)
     OR ROM64_INSTR_PT(31) OR ROM64_INSTR_PT(38)
     OR ROM64_INSTR_PT(41) OR ROM64_INSTR_PT(49)
     OR ROM64_INSTR_PT(51) OR ROM64_INSTR_PT(52)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(61)
     OR ROM64_INSTR_PT(64) OR ROM64_INSTR_PT(70)
     OR ROM64_INSTR_PT(71) OR ROM64_INSTR_PT(75)
     OR ROM64_INSTR_PT(76) OR ROM64_INSTR_PT(83)
     OR ROM64_INSTR_PT(86) OR ROM64_INSTR_PT(90)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(97)
     OR ROM64_INSTR_PT(99) OR ROM64_INSTR_PT(100)
     OR ROM64_INSTR_PT(102) OR ROM64_INSTR_PT(105)
     OR ROM64_INSTR_PT(113) OR ROM64_INSTR_PT(115)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(124) OR ROM64_INSTR_PT(127)
     OR ROM64_INSTR_PT(132) OR ROM64_INSTR_PT(133)
     OR ROM64_INSTR_PT(134) OR ROM64_INSTR_PT(136)
     OR ROM64_INSTR_PT(137) OR ROM64_INSTR_PT(140)
     OR ROM64_INSTR_PT(144) OR ROM64_INSTR_PT(148)
     OR ROM64_INSTR_PT(153) OR ROM64_INSTR_PT(158)
     OR ROM64_INSTR_PT(164) OR ROM64_INSTR_PT(168)
     OR ROM64_INSTR_PT(169) OR ROM64_INSTR_PT(171)
     OR ROM64_INSTR_PT(172) OR ROM64_INSTR_PT(181)
     OR ROM64_INSTR_PT(184) OR ROM64_INSTR_PT(185)
     OR ROM64_INSTR_PT(186) OR ROM64_INSTR_PT(194)
     OR ROM64_INSTR_PT(199) OR ROM64_INSTR_PT(202)
     OR ROM64_INSTR_PT(204) OR ROM64_INSTR_PT(211)
     OR ROM64_INSTR_PT(215) OR ROM64_INSTR_PT(217)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(219)
     OR ROM64_INSTR_PT(222) OR ROM64_INSTR_PT(226)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(238) OR ROM64_INSTR_PT(241)
     OR ROM64_INSTR_PT(245) OR ROM64_INSTR_PT(252)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(263) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(270)
     OR ROM64_INSTR_PT(271) OR ROM64_INSTR_PT(272)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(275)
     OR ROM64_INSTR_PT(276) OR ROM64_INSTR_PT(277)
     OR ROM64_INSTR_PT(282) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(285) OR ROM64_INSTR_PT(287)
     OR ROM64_INSTR_PT(293) OR ROM64_INSTR_PT(294)
     OR ROM64_INSTR_PT(297) OR ROM64_INSTR_PT(298)
     OR ROM64_INSTR_PT(299) OR ROM64_INSTR_PT(302)
     OR ROM64_INSTR_PT(305) OR ROM64_INSTR_PT(308)
     OR ROM64_INSTR_PT(311) OR ROM64_INSTR_PT(312)
     OR ROM64_INSTR_PT(315) OR ROM64_INSTR_PT(319)
     OR ROM64_INSTR_PT(324) OR ROM64_INSTR_PT(325)
     OR ROM64_INSTR_PT(331) OR ROM64_INSTR_PT(340)
     OR ROM64_INSTR_PT(361) OR ROM64_INSTR_PT(364)
     OR ROM64_INSTR_PT(374) OR ROM64_INSTR_PT(375)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(383)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(385)
     OR ROM64_INSTR_PT(388) OR ROM64_INSTR_PT(391)
     OR ROM64_INSTR_PT(394) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(403) OR ROM64_INSTR_PT(404)
     OR ROM64_INSTR_PT(406) OR ROM64_INSTR_PT(410)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(424) OR ROM64_INSTR_PT(428)
     OR ROM64_INSTR_PT(430) OR ROM64_INSTR_PT(432)
     OR ROM64_INSTR_PT(434) OR ROM64_INSTR_PT(437)
     OR ROM64_INSTR_PT(438) OR ROM64_INSTR_PT(439)
     OR ROM64_INSTR_PT(440) OR ROM64_INSTR_PT(441)
     OR ROM64_INSTR_PT(443) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(453)
     OR ROM64_INSTR_PT(454) OR ROM64_INSTR_PT(455)
     OR ROM64_INSTR_PT(468) OR ROM64_INSTR_PT(478)
     OR ROM64_INSTR_PT(481) OR ROM64_INSTR_PT(482)
     OR ROM64_INSTR_PT(484) OR ROM64_INSTR_PT(485)
     OR ROM64_INSTR_PT(493) OR ROM64_INSTR_PT(495)
     OR ROM64_INSTR_PT(496) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(505)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(510)
     OR ROM64_INSTR_PT(511) OR ROM64_INSTR_PT(512)
     OR ROM64_INSTR_PT(516) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(521) OR ROM64_INSTR_PT(522)
     OR ROM64_INSTR_PT(525) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(531) OR ROM64_INSTR_PT(532)
     OR ROM64_INSTR_PT(534) OR ROM64_INSTR_PT(535)
     OR ROM64_INSTR_PT(544) OR ROM64_INSTR_PT(545)
     OR ROM64_INSTR_PT(546) OR ROM64_INSTR_PT(549)
     OR ROM64_INSTR_PT(552) OR ROM64_INSTR_PT(555)
     OR ROM64_INSTR_PT(558) OR ROM64_INSTR_PT(559)
     OR ROM64_INSTR_PT(563) OR ROM64_INSTR_PT(564)
     OR ROM64_INSTR_PT(566) OR ROM64_INSTR_PT(569)
     OR ROM64_INSTR_PT(571) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(581)
     OR ROM64_INSTR_PT(582) OR ROM64_INSTR_PT(583)
     OR ROM64_INSTR_PT(586) OR ROM64_INSTR_PT(587)
     OR ROM64_INSTR_PT(588) OR ROM64_INSTR_PT(589)
     OR ROM64_INSTR_PT(591) OR ROM64_INSTR_PT(595)
     OR ROM64_INSTR_PT(600) OR ROM64_INSTR_PT(604)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(607)
     OR ROM64_INSTR_PT(608) OR ROM64_INSTR_PT(615)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(625)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(629) OR ROM64_INSTR_PT(632)
     OR ROM64_INSTR_PT(633) OR ROM64_INSTR_PT(639)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(644)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(664)
     OR ROM64_INSTR_PT(666) OR ROM64_INSTR_PT(678)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(698)
     OR ROM64_INSTR_PT(702) OR ROM64_INSTR_PT(722)
     OR ROM64_INSTR_PT(728) OR ROM64_INSTR_PT(731)
     OR ROM64_INSTR_PT(735) OR ROM64_INSTR_PT(738)
     OR ROM64_INSTR_PT(744) OR ROM64_INSTR_PT(761)
     OR ROM64_INSTR_PT(769) OR ROM64_INSTR_PT(776)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(832)
     OR ROM64_INSTR_PT(846) OR ROM64_INSTR_PT(854)
     OR ROM64_INSTR_PT(856) OR ROM64_INSTR_PT(864)
     OR ROM64_INSTR_PT(870));
MQQ921:TEMPLATE(30) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(7) OR ROM64_INSTR_PT(9)
     OR ROM64_INSTR_PT(10) OR ROM64_INSTR_PT(14)
     OR ROM64_INSTR_PT(17) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(38) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(50)
     OR ROM64_INSTR_PT(51) OR ROM64_INSTR_PT(52)
     OR ROM64_INSTR_PT(55) OR ROM64_INSTR_PT(61)
     OR ROM64_INSTR_PT(64) OR ROM64_INSTR_PT(70)
     OR ROM64_INSTR_PT(71) OR ROM64_INSTR_PT(75)
     OR ROM64_INSTR_PT(76) OR ROM64_INSTR_PT(77)
     OR ROM64_INSTR_PT(78) OR ROM64_INSTR_PT(80)
     OR ROM64_INSTR_PT(83) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(86) OR ROM64_INSTR_PT(89)
     OR ROM64_INSTR_PT(90) OR ROM64_INSTR_PT(92)
     OR ROM64_INSTR_PT(96) OR ROM64_INSTR_PT(99)
     OR ROM64_INSTR_PT(100) OR ROM64_INSTR_PT(102)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(105)
     OR ROM64_INSTR_PT(106) OR ROM64_INSTR_PT(110)
     OR ROM64_INSTR_PT(113) OR ROM64_INSTR_PT(114)
     OR ROM64_INSTR_PT(115) OR ROM64_INSTR_PT(116)
     OR ROM64_INSTR_PT(117) OR ROM64_INSTR_PT(118)
     OR ROM64_INSTR_PT(121) OR ROM64_INSTR_PT(124)
     OR ROM64_INSTR_PT(127) OR ROM64_INSTR_PT(132)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(143)
     OR ROM64_INSTR_PT(144) OR ROM64_INSTR_PT(148)
     OR ROM64_INSTR_PT(153) OR ROM64_INSTR_PT(169)
     OR ROM64_INSTR_PT(171) OR ROM64_INSTR_PT(175)
     OR ROM64_INSTR_PT(177) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(181) OR ROM64_INSTR_PT(183)
     OR ROM64_INSTR_PT(184) OR ROM64_INSTR_PT(185)
     OR ROM64_INSTR_PT(186) OR ROM64_INSTR_PT(188)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(199)
     OR ROM64_INSTR_PT(202) OR ROM64_INSTR_PT(204)
     OR ROM64_INSTR_PT(208) OR ROM64_INSTR_PT(213)
     OR ROM64_INSTR_PT(214) OR ROM64_INSTR_PT(215)
     OR ROM64_INSTR_PT(217) OR ROM64_INSTR_PT(218)
     OR ROM64_INSTR_PT(221) OR ROM64_INSTR_PT(222)
     OR ROM64_INSTR_PT(223) OR ROM64_INSTR_PT(226)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(233) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(241) OR ROM64_INSTR_PT(252)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(263) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(270)
     OR ROM64_INSTR_PT(271) OR ROM64_INSTR_PT(274)
     OR ROM64_INSTR_PT(275) OR ROM64_INSTR_PT(276)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(282)
     OR ROM64_INSTR_PT(285) OR ROM64_INSTR_PT(286)
     OR ROM64_INSTR_PT(293) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(298) OR ROM64_INSTR_PT(299)
     OR ROM64_INSTR_PT(302) OR ROM64_INSTR_PT(305)
     OR ROM64_INSTR_PT(308) OR ROM64_INSTR_PT(315)
     OR ROM64_INSTR_PT(319) OR ROM64_INSTR_PT(322)
     OR ROM64_INSTR_PT(331) OR ROM64_INSTR_PT(339)
     OR ROM64_INSTR_PT(347) OR ROM64_INSTR_PT(349)
     OR ROM64_INSTR_PT(350) OR ROM64_INSTR_PT(358)
     OR ROM64_INSTR_PT(364) OR ROM64_INSTR_PT(367)
     OR ROM64_INSTR_PT(369) OR ROM64_INSTR_PT(371)
     OR ROM64_INSTR_PT(374) OR ROM64_INSTR_PT(375)
     OR ROM64_INSTR_PT(378) OR ROM64_INSTR_PT(379)
     OR ROM64_INSTR_PT(383) OR ROM64_INSTR_PT(385)
     OR ROM64_INSTR_PT(391) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(397) OR ROM64_INSTR_PT(403)
     OR ROM64_INSTR_PT(404) OR ROM64_INSTR_PT(410)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(424)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(432) OR ROM64_INSTR_PT(434)
     OR ROM64_INSTR_PT(435) OR ROM64_INSTR_PT(437)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(453)
     OR ROM64_INSTR_PT(461) OR ROM64_INSTR_PT(463)
     OR ROM64_INSTR_PT(466) OR ROM64_INSTR_PT(478)
     OR ROM64_INSTR_PT(481) OR ROM64_INSTR_PT(482)
     OR ROM64_INSTR_PT(484) OR ROM64_INSTR_PT(485)
     OR ROM64_INSTR_PT(493) OR ROM64_INSTR_PT(495)
     OR ROM64_INSTR_PT(496) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(505)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(510)
     OR ROM64_INSTR_PT(511) OR ROM64_INSTR_PT(512)
     OR ROM64_INSTR_PT(521) OR ROM64_INSTR_PT(522)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(525)
     OR ROM64_INSTR_PT(534) OR ROM64_INSTR_PT(540)
     OR ROM64_INSTR_PT(545) OR ROM64_INSTR_PT(546)
     OR ROM64_INSTR_PT(552) OR ROM64_INSTR_PT(555)
     OR ROM64_INSTR_PT(557) OR ROM64_INSTR_PT(558)
     OR ROM64_INSTR_PT(559) OR ROM64_INSTR_PT(563)
     OR ROM64_INSTR_PT(569) OR ROM64_INSTR_PT(571)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(582) OR ROM64_INSTR_PT(583)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(588)
     OR ROM64_INSTR_PT(591) OR ROM64_INSTR_PT(592)
     OR ROM64_INSTR_PT(595) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(600) OR ROM64_INSTR_PT(606)
     OR ROM64_INSTR_PT(608) OR ROM64_INSTR_PT(609)
     OR ROM64_INSTR_PT(613) OR ROM64_INSTR_PT(615)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(619)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(629)
     OR ROM64_INSTR_PT(632) OR ROM64_INSTR_PT(633)
     OR ROM64_INSTR_PT(639) OR ROM64_INSTR_PT(642)
     OR ROM64_INSTR_PT(644) OR ROM64_INSTR_PT(666)
     OR ROM64_INSTR_PT(678) OR ROM64_INSTR_PT(685)
     OR ROM64_INSTR_PT(687) OR ROM64_INSTR_PT(691)
     OR ROM64_INSTR_PT(695) OR ROM64_INSTR_PT(716)
     OR ROM64_INSTR_PT(722) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(728)
     OR ROM64_INSTR_PT(731) OR ROM64_INSTR_PT(733)
     OR ROM64_INSTR_PT(735) OR ROM64_INSTR_PT(736)
     OR ROM64_INSTR_PT(738) OR ROM64_INSTR_PT(744)
     OR ROM64_INSTR_PT(761) OR ROM64_INSTR_PT(769)
     OR ROM64_INSTR_PT(770) OR ROM64_INSTR_PT(776)
     OR ROM64_INSTR_PT(834) OR ROM64_INSTR_PT(846)
     OR ROM64_INSTR_PT(856) OR ROM64_INSTR_PT(864)
     OR ROM64_INSTR_PT(870));
MQQ922:TEMPLATE(31) <= 
    (ROM64_INSTR_PT(33) OR ROM64_INSTR_PT(60)
     OR ROM64_INSTR_PT(79) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(103) OR ROM64_INSTR_PT(142)
     OR ROM64_INSTR_PT(147) OR ROM64_INSTR_PT(150)
     OR ROM64_INSTR_PT(160) OR ROM64_INSTR_PT(168)
     OR ROM64_INSTR_PT(176) OR ROM64_INSTR_PT(187)
     OR ROM64_INSTR_PT(207) OR ROM64_INSTR_PT(209)
     OR ROM64_INSTR_PT(219) OR ROM64_INSTR_PT(224)
     OR ROM64_INSTR_PT(228) OR ROM64_INSTR_PT(231)
     OR ROM64_INSTR_PT(247) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(281) OR ROM64_INSTR_PT(288)
     OR ROM64_INSTR_PT(296) OR ROM64_INSTR_PT(304)
     OR ROM64_INSTR_PT(309) OR ROM64_INSTR_PT(314)
     OR ROM64_INSTR_PT(327) OR ROM64_INSTR_PT(332)
     OR ROM64_INSTR_PT(341) OR ROM64_INSTR_PT(352)
     OR ROM64_INSTR_PT(361) OR ROM64_INSTR_PT(374)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(406)
     OR ROM64_INSTR_PT(464) OR ROM64_INSTR_PT(471)
     OR ROM64_INSTR_PT(491) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(632) OR ROM64_INSTR_PT(635)
     OR ROM64_INSTR_PT(641) OR ROM64_INSTR_PT(654)
     OR ROM64_INSTR_PT(675) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(728)
     OR ROM64_INSTR_PT(733) OR ROM64_INSTR_PT(735)
     OR ROM64_INSTR_PT(738) OR ROM64_INSTR_PT(759)
     OR ROM64_INSTR_PT(766) OR ROM64_INSTR_PT(781)
     OR ROM64_INSTR_PT(794) OR ROM64_INSTR_PT(809)
    );
MQQ923:UCODE_END <= 
    (ROM64_INSTR_PT(198) OR ROM64_INSTR_PT(200)
     OR ROM64_INSTR_PT(212) OR ROM64_INSTR_PT(386)
     OR ROM64_INSTR_PT(443) OR ROM64_INSTR_PT(444)
     OR ROM64_INSTR_PT(452) OR ROM64_INSTR_PT(516)
     OR ROM64_INSTR_PT(518) OR ROM64_INSTR_PT(528)
     OR ROM64_INSTR_PT(542) OR ROM64_INSTR_PT(550)
     OR ROM64_INSTR_PT(556) OR ROM64_INSTR_PT(560)
     OR ROM64_INSTR_PT(567) OR ROM64_INSTR_PT(574)
     OR ROM64_INSTR_PT(577) OR ROM64_INSTR_PT(578)
     OR ROM64_INSTR_PT(581) OR ROM64_INSTR_PT(593)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(606)
     OR ROM64_INSTR_PT(607) OR ROM64_INSTR_PT(622)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(668)
     OR ROM64_INSTR_PT(690) OR ROM64_INSTR_PT(699)
     OR ROM64_INSTR_PT(704) OR ROM64_INSTR_PT(706)
     OR ROM64_INSTR_PT(714) OR ROM64_INSTR_PT(718)
     OR ROM64_INSTR_PT(741) OR ROM64_INSTR_PT(785)
     OR ROM64_INSTR_PT(790) OR ROM64_INSTR_PT(813)
     OR ROM64_INSTR_PT(823) OR ROM64_INSTR_PT(824)
     OR ROM64_INSTR_PT(826) OR ROM64_INSTR_PT(828)
     OR ROM64_INSTR_PT(841) OR ROM64_INSTR_PT(844)
     OR ROM64_INSTR_PT(845) OR ROM64_INSTR_PT(849)
     OR ROM64_INSTR_PT(854));
MQQ924:UCODE_END_EARLY <= 
    (ROM64_INSTR_PT(376) OR ROM64_INSTR_PT(390)
     OR ROM64_INSTR_PT(650) OR ROM64_INSTR_PT(676)
     OR ROM64_INSTR_PT(683) OR ROM64_INSTR_PT(689)
     OR ROM64_INSTR_PT(730) OR ROM64_INSTR_PT(742)
     OR ROM64_INSTR_PT(757) OR ROM64_INSTR_PT(760)
     OR ROM64_INSTR_PT(787) OR ROM64_INSTR_PT(788)
     OR ROM64_INSTR_PT(800) OR ROM64_INSTR_PT(802)
     OR ROM64_INSTR_PT(803) OR ROM64_INSTR_PT(807)
     OR ROM64_INSTR_PT(814) OR ROM64_INSTR_PT(818)
     OR ROM64_INSTR_PT(825) OR ROM64_INSTR_PT(830)
     OR ROM64_INSTR_PT(874));
MQQ925:LOOP_BEGIN <= 
    (ROM64_INSTR_PT(26) OR ROM64_INSTR_PT(55)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(124)
     OR ROM64_INSTR_PT(147) OR ROM64_INSTR_PT(210)
     OR ROM64_INSTR_PT(228) OR ROM64_INSTR_PT(231)
     OR ROM64_INSTR_PT(239) OR ROM64_INSTR_PT(246)
     OR ROM64_INSTR_PT(255) OR ROM64_INSTR_PT(306)
     OR ROM64_INSTR_PT(310) OR ROM64_INSTR_PT(316)
     OR ROM64_INSTR_PT(322) OR ROM64_INSTR_PT(349)
     OR ROM64_INSTR_PT(369) OR ROM64_INSTR_PT(379)
     OR ROM64_INSTR_PT(411) OR ROM64_INSTR_PT(412)
     OR ROM64_INSTR_PT(436) OR ROM64_INSTR_PT(450)
     OR ROM64_INSTR_PT(462) OR ROM64_INSTR_PT(487)
     OR ROM64_INSTR_PT(493) OR ROM64_INSTR_PT(496)
     OR ROM64_INSTR_PT(546) OR ROM64_INSTR_PT(559)
     OR ROM64_INSTR_PT(572) OR ROM64_INSTR_PT(590)
     OR ROM64_INSTR_PT(610));
MQQ926:LOOP_END <= 
    (ROM64_INSTR_PT(149) OR ROM64_INSTR_PT(156)
     OR ROM64_INSTR_PT(376) OR ROM64_INSTR_PT(469)
     OR ROM64_INSTR_PT(494) OR ROM64_INSTR_PT(502)
     OR ROM64_INSTR_PT(565) OR ROM64_INSTR_PT(638)
     OR ROM64_INSTR_PT(647) OR ROM64_INSTR_PT(656)
     OR ROM64_INSTR_PT(680) OR ROM64_INSTR_PT(701)
     OR ROM64_INSTR_PT(751) OR ROM64_INSTR_PT(775)
     OR ROM64_INSTR_PT(779) OR ROM64_INSTR_PT(789)
     OR ROM64_INSTR_PT(799) OR ROM64_INSTR_PT(807)
     OR ROM64_INSTR_PT(815) OR ROM64_INSTR_PT(816)
     OR ROM64_INSTR_PT(850) OR ROM64_INSTR_PT(862)
     OR ROM64_INSTR_PT(875));
MQQ927:COUNT_SRC(0) <= 
    (ROM64_INSTR_PT(72) OR ROM64_INSTR_PT(752)
     OR ROM64_INSTR_PT(768) OR ROM64_INSTR_PT(876)
     OR ROM64_INSTR_PT(881) OR ROM64_INSTR_PT(882)
     OR ROM64_INSTR_PT(887) OR ROM64_INSTR_PT(888)
     OR ROM64_INSTR_PT(889));
MQQ928:COUNT_SRC(1) <= 
    (ROM64_INSTR_PT(839) OR ROM64_INSTR_PT(879)
     OR ROM64_INSTR_PT(882) OR ROM64_INSTR_PT(884)
     OR ROM64_INSTR_PT(885) OR ROM64_INSTR_PT(888)
     OR ROM64_INSTR_PT(889));
MQQ929:COUNT_SRC(2) <= 
    (ROM64_INSTR_PT(686) OR ROM64_INSTR_PT(752)
     OR ROM64_INSTR_PT(768) OR ROM64_INSTR_PT(831)
     OR ROM64_INSTR_PT(839) OR ROM64_INSTR_PT(887)
     OR ROM64_INSTR_PT(888) OR ROM64_INSTR_PT(889)
    );
MQQ930:EXTRT <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(6)
     OR ROM64_INSTR_PT(19) OR ROM64_INSTR_PT(24)
     OR ROM64_INSTR_PT(27) OR ROM64_INSTR_PT(47)
     OR ROM64_INSTR_PT(48) OR ROM64_INSTR_PT(63)
     OR ROM64_INSTR_PT(69) OR ROM64_INSTR_PT(74)
     OR ROM64_INSTR_PT(91) OR ROM64_INSTR_PT(95)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(107)
     OR ROM64_INSTR_PT(120) OR ROM64_INSTR_PT(123)
     OR ROM64_INSTR_PT(130) OR ROM64_INSTR_PT(131)
     OR ROM64_INSTR_PT(133) OR ROM64_INSTR_PT(135)
     OR ROM64_INSTR_PT(138) OR ROM64_INSTR_PT(140)
     OR ROM64_INSTR_PT(141) OR ROM64_INSTR_PT(151)
     OR ROM64_INSTR_PT(152) OR ROM64_INSTR_PT(159)
     OR ROM64_INSTR_PT(163) OR ROM64_INSTR_PT(164)
     OR ROM64_INSTR_PT(167) OR ROM64_INSTR_PT(189)
     OR ROM64_INSTR_PT(192) OR ROM64_INSTR_PT(220)
     OR ROM64_INSTR_PT(227) OR ROM64_INSTR_PT(234)
     OR ROM64_INSTR_PT(235) OR ROM64_INSTR_PT(250)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(258)
     OR ROM64_INSTR_PT(266) OR ROM64_INSTR_PT(267)
     OR ROM64_INSTR_PT(279) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(300) OR ROM64_INSTR_PT(301)
     OR ROM64_INSTR_PT(303) OR ROM64_INSTR_PT(317)
     OR ROM64_INSTR_PT(318) OR ROM64_INSTR_PT(328)
     OR ROM64_INSTR_PT(330) OR ROM64_INSTR_PT(331)
     OR ROM64_INSTR_PT(335) OR ROM64_INSTR_PT(337)
     OR ROM64_INSTR_PT(338) OR ROM64_INSTR_PT(344)
     OR ROM64_INSTR_PT(355) OR ROM64_INSTR_PT(356)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(393)
     OR ROM64_INSTR_PT(394) OR ROM64_INSTR_PT(398)
     OR ROM64_INSTR_PT(418) OR ROM64_INSTR_PT(423)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(447)
     OR ROM64_INSTR_PT(449) OR ROM64_INSTR_PT(476)
     OR ROM64_INSTR_PT(486) OR ROM64_INSTR_PT(487)
     OR ROM64_INSTR_PT(496) OR ROM64_INSTR_PT(500)
     OR ROM64_INSTR_PT(501) OR ROM64_INSTR_PT(526)
     OR ROM64_INSTR_PT(547) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(594) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(624) OR ROM64_INSTR_PT(630)
     OR ROM64_INSTR_PT(631) OR ROM64_INSTR_PT(640)
     OR ROM64_INSTR_PT(651) OR ROM64_INSTR_PT(665)
     OR ROM64_INSTR_PT(670) OR ROM64_INSTR_PT(671)
     OR ROM64_INSTR_PT(672) OR ROM64_INSTR_PT(673)
     OR ROM64_INSTR_PT(674) OR ROM64_INSTR_PT(688)
     OR ROM64_INSTR_PT(696) OR ROM64_INSTR_PT(700)
     OR ROM64_INSTR_PT(707) OR ROM64_INSTR_PT(712)
     OR ROM64_INSTR_PT(727) OR ROM64_INSTR_PT(732)
     OR ROM64_INSTR_PT(737) OR ROM64_INSTR_PT(743)
     OR ROM64_INSTR_PT(744) OR ROM64_INSTR_PT(746)
     OR ROM64_INSTR_PT(747) OR ROM64_INSTR_PT(750)
     OR ROM64_INSTR_PT(755) OR ROM64_INSTR_PT(756)
     OR ROM64_INSTR_PT(763) OR ROM64_INSTR_PT(764)
     OR ROM64_INSTR_PT(767) OR ROM64_INSTR_PT(771)
     OR ROM64_INSTR_PT(774) OR ROM64_INSTR_PT(776)
     OR ROM64_INSTR_PT(777) OR ROM64_INSTR_PT(780)
     OR ROM64_INSTR_PT(782) OR ROM64_INSTR_PT(783)
     OR ROM64_INSTR_PT(784) OR ROM64_INSTR_PT(786)
     OR ROM64_INSTR_PT(793) OR ROM64_INSTR_PT(795)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(810)
     OR ROM64_INSTR_PT(812) OR ROM64_INSTR_PT(820)
     OR ROM64_INSTR_PT(821) OR ROM64_INSTR_PT(833)
     OR ROM64_INSTR_PT(835) OR ROM64_INSTR_PT(837)
     OR ROM64_INSTR_PT(838) OR ROM64_INSTR_PT(848)
     OR ROM64_INSTR_PT(857) OR ROM64_INSTR_PT(859)
     OR ROM64_INSTR_PT(860) OR ROM64_INSTR_PT(863)
     OR ROM64_INSTR_PT(864) OR ROM64_INSTR_PT(865)
     OR ROM64_INSTR_PT(866) OR ROM64_INSTR_PT(867)
     OR ROM64_INSTR_PT(868) OR ROM64_INSTR_PT(871)
     OR ROM64_INSTR_PT(877) OR ROM64_INSTR_PT(878)
     OR ROM64_INSTR_PT(880));
MQQ931:EXTS1 <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(19)
     OR ROM64_INSTR_PT(32) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(47) OR ROM64_INSTR_PT(74)
     OR ROM64_INSTR_PT(81) OR ROM64_INSTR_PT(91)
     OR ROM64_INSTR_PT(94) OR ROM64_INSTR_PT(100)
     OR ROM64_INSTR_PT(131) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(138) OR ROM64_INSTR_PT(159)
     OR ROM64_INSTR_PT(165) OR ROM64_INSTR_PT(167)
     OR ROM64_INSTR_PT(193) OR ROM64_INSTR_PT(211)
     OR ROM64_INSTR_PT(225) OR ROM64_INSTR_PT(227)
     OR ROM64_INSTR_PT(232) OR ROM64_INSTR_PT(235)
     OR ROM64_INSTR_PT(279) OR ROM64_INSTR_PT(289)
     OR ROM64_INSTR_PT(291) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(300) OR ROM64_INSTR_PT(301)
     OR ROM64_INSTR_PT(317) OR ROM64_INSTR_PT(318)
     OR ROM64_INSTR_PT(326) OR ROM64_INSTR_PT(328)
     OR ROM64_INSTR_PT(330) OR ROM64_INSTR_PT(331)
     OR ROM64_INSTR_PT(335) OR ROM64_INSTR_PT(337)
     OR ROM64_INSTR_PT(338) OR ROM64_INSTR_PT(344)
     OR ROM64_INSTR_PT(350) OR ROM64_INSTR_PT(358)
     OR ROM64_INSTR_PT(373) OR ROM64_INSTR_PT(379)
     OR ROM64_INSTR_PT(393) OR ROM64_INSTR_PT(398)
     OR ROM64_INSTR_PT(400) OR ROM64_INSTR_PT(421)
     OR ROM64_INSTR_PT(438) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(449) OR ROM64_INSTR_PT(465)
     OR ROM64_INSTR_PT(476) OR ROM64_INSTR_PT(479)
     OR ROM64_INSTR_PT(486) OR ROM64_INSTR_PT(500)
     OR ROM64_INSTR_PT(526) OR ROM64_INSTR_PT(543)
     OR ROM64_INSTR_PT(566) OR ROM64_INSTR_PT(577)
     OR ROM64_INSTR_PT(581) OR ROM64_INSTR_PT(593)
     OR ROM64_INSTR_PT(594) OR ROM64_INSTR_PT(604)
     OR ROM64_INSTR_PT(624) OR ROM64_INSTR_PT(630)
     OR ROM64_INSTR_PT(631) OR ROM64_INSTR_PT(652)
     OR ROM64_INSTR_PT(669) OR ROM64_INSTR_PT(671)
     OR ROM64_INSTR_PT(672) OR ROM64_INSTR_PT(673)
     OR ROM64_INSTR_PT(674) OR ROM64_INSTR_PT(688)
     OR ROM64_INSTR_PT(692) OR ROM64_INSTR_PT(694)
     OR ROM64_INSTR_PT(697) OR ROM64_INSTR_PT(700)
     OR ROM64_INSTR_PT(707) OR ROM64_INSTR_PT(708)
     OR ROM64_INSTR_PT(710) OR ROM64_INSTR_PT(712)
     OR ROM64_INSTR_PT(715) OR ROM64_INSTR_PT(720)
     OR ROM64_INSTR_PT(725) OR ROM64_INSTR_PT(732)
     OR ROM64_INSTR_PT(737) OR ROM64_INSTR_PT(741)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(746)
     OR ROM64_INSTR_PT(747) OR ROM64_INSTR_PT(749)
     OR ROM64_INSTR_PT(750) OR ROM64_INSTR_PT(755)
     OR ROM64_INSTR_PT(758) OR ROM64_INSTR_PT(762)
     OR ROM64_INSTR_PT(763) OR ROM64_INSTR_PT(764)
     OR ROM64_INSTR_PT(767) OR ROM64_INSTR_PT(771)
     OR ROM64_INSTR_PT(774) OR ROM64_INSTR_PT(777)
     OR ROM64_INSTR_PT(778) OR ROM64_INSTR_PT(780)
     OR ROM64_INSTR_PT(782) OR ROM64_INSTR_PT(783)
     OR ROM64_INSTR_PT(784) OR ROM64_INSTR_PT(786)
     OR ROM64_INSTR_PT(793) OR ROM64_INSTR_PT(795)
     OR ROM64_INSTR_PT(796) OR ROM64_INSTR_PT(806)
     OR ROM64_INSTR_PT(810) OR ROM64_INSTR_PT(812)
     OR ROM64_INSTR_PT(817) OR ROM64_INSTR_PT(820)
     OR ROM64_INSTR_PT(821) OR ROM64_INSTR_PT(823)
     OR ROM64_INSTR_PT(828) OR ROM64_INSTR_PT(835)
     OR ROM64_INSTR_PT(836) OR ROM64_INSTR_PT(837)
     OR ROM64_INSTR_PT(838) OR ROM64_INSTR_PT(842)
     OR ROM64_INSTR_PT(843) OR ROM64_INSTR_PT(844)
     OR ROM64_INSTR_PT(847) OR ROM64_INSTR_PT(848)
     OR ROM64_INSTR_PT(849) OR ROM64_INSTR_PT(851)
     OR ROM64_INSTR_PT(853) OR ROM64_INSTR_PT(859)
     OR ROM64_INSTR_PT(861) OR ROM64_INSTR_PT(865)
     OR ROM64_INSTR_PT(866) OR ROM64_INSTR_PT(867)
     OR ROM64_INSTR_PT(871) OR ROM64_INSTR_PT(877)
     OR ROM64_INSTR_PT(880));
MQQ932:EXTS2 <= 
    (ROM64_INSTR_PT(23) OR ROM64_INSTR_PT(27)
     OR ROM64_INSTR_PT(44) OR ROM64_INSTR_PT(47)
     OR ROM64_INSTR_PT(88) OR ROM64_INSTR_PT(91)
     OR ROM64_INSTR_PT(131) OR ROM64_INSTR_PT(138)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(152)
     OR ROM64_INSTR_PT(167) OR ROM64_INSTR_PT(178)
     OR ROM64_INSTR_PT(182) OR ROM64_INSTR_PT(189)
     OR ROM64_INSTR_PT(211) OR ROM64_INSTR_PT(298)
     OR ROM64_INSTR_PT(318) OR ROM64_INSTR_PT(330)
     OR ROM64_INSTR_PT(331) OR ROM64_INSTR_PT(335)
     OR ROM64_INSTR_PT(337) OR ROM64_INSTR_PT(344)
     OR ROM64_INSTR_PT(346) OR ROM64_INSTR_PT(350)
     OR ROM64_INSTR_PT(356) OR ROM64_INSTR_PT(358)
     OR ROM64_INSTR_PT(373) OR ROM64_INSTR_PT(380)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(400) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(432) OR ROM64_INSTR_PT(441)
     OR ROM64_INSTR_PT(479) OR ROM64_INSTR_PT(500)
     OR ROM64_INSTR_PT(516) OR ROM64_INSTR_PT(526)
     OR ROM64_INSTR_PT(530) OR ROM64_INSTR_PT(542)
     OR ROM64_INSTR_PT(577) OR ROM64_INSTR_PT(580)
     OR ROM64_INSTR_PT(581) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(627)
     OR ROM64_INSTR_PT(631) OR ROM64_INSTR_PT(652)
     OR ROM64_INSTR_PT(672) OR ROM64_INSTR_PT(674)
     OR ROM64_INSTR_PT(696) OR ROM64_INSTR_PT(697)
     OR ROM64_INSTR_PT(700) OR ROM64_INSTR_PT(707)
     OR ROM64_INSTR_PT(715) OR ROM64_INSTR_PT(718)
     OR ROM64_INSTR_PT(725) OR ROM64_INSTR_PT(737)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(744)
     OR ROM64_INSTR_PT(745) OR ROM64_INSTR_PT(746)
     OR ROM64_INSTR_PT(750) OR ROM64_INSTR_PT(754)
     OR ROM64_INSTR_PT(756) OR ROM64_INSTR_PT(758)
     OR ROM64_INSTR_PT(763) OR ROM64_INSTR_PT(765)
     OR ROM64_INSTR_PT(767) OR ROM64_INSTR_PT(771)
     OR ROM64_INSTR_PT(772) OR ROM64_INSTR_PT(774)
     OR ROM64_INSTR_PT(776) OR ROM64_INSTR_PT(778)
     OR ROM64_INSTR_PT(784) OR ROM64_INSTR_PT(786)
     OR ROM64_INSTR_PT(812) OR ROM64_INSTR_PT(813)
     OR ROM64_INSTR_PT(820) OR ROM64_INSTR_PT(823)
     OR ROM64_INSTR_PT(828) OR ROM64_INSTR_PT(842)
     OR ROM64_INSTR_PT(843) OR ROM64_INSTR_PT(848)
     OR ROM64_INSTR_PT(854) OR ROM64_INSTR_PT(859)
     OR ROM64_INSTR_PT(860) OR ROM64_INSTR_PT(863)
     OR ROM64_INSTR_PT(866) OR ROM64_INSTR_PT(867)
     OR ROM64_INSTR_PT(868) OR ROM64_INSTR_PT(877)
     OR ROM64_INSTR_PT(880));
MQQ933:EXTS3 <= 
    (ROM64_INSTR_PT(47) OR ROM64_INSTR_PT(94)
     OR ROM64_INSTR_PT(100) OR ROM64_INSTR_PT(135)
     OR ROM64_INSTR_PT(159) OR ROM64_INSTR_PT(163)
     OR ROM64_INSTR_PT(192) OR ROM64_INSTR_PT(225)
     OR ROM64_INSTR_PT(235) OR ROM64_INSTR_PT(251)
     OR ROM64_INSTR_PT(279) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(300) OR ROM64_INSTR_PT(326)
     OR ROM64_INSTR_PT(337) OR ROM64_INSTR_PT(338)
     OR ROM64_INSTR_PT(350) OR ROM64_INSTR_PT(358)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(384)
     OR ROM64_INSTR_PT(398) OR ROM64_INSTR_PT(413)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(447)
     OR ROM64_INSTR_PT(524) OR ROM64_INSTR_PT(526)
     OR ROM64_INSTR_PT(561) OR ROM64_INSTR_PT(572)
     OR ROM64_INSTR_PT(594) OR ROM64_INSTR_PT(630)
     OR ROM64_INSTR_PT(670) OR ROM64_INSTR_PT(692)
     OR ROM64_INSTR_PT(697) OR ROM64_INSTR_PT(712)
     OR ROM64_INSTR_PT(715) OR ROM64_INSTR_PT(749)
     OR ROM64_INSTR_PT(758) OR ROM64_INSTR_PT(778)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(833)
     OR ROM64_INSTR_PT(837) OR ROM64_INSTR_PT(838)
     OR ROM64_INSTR_PT(871));
MQQ934:SEL0_5 <= 
    (ROM64_INSTR_PT(652) OR ROM64_INSTR_PT(718)
    );
MQQ935:SEL6_10(0) <= 
    (ROM64_INSTR_PT(40) OR ROM64_INSTR_PT(69)
     OR ROM64_INSTR_PT(82) OR ROM64_INSTR_PT(95)
     OR ROM64_INSTR_PT(107) OR ROM64_INSTR_PT(200)
     OR ROM64_INSTR_PT(211) OR ROM64_INSTR_PT(267)
     OR ROM64_INSTR_PT(386) OR ROM64_INSTR_PT(443)
     OR ROM64_INSTR_PT(444) OR ROM64_INSTR_PT(452)
     OR ROM64_INSTR_PT(516) OR ROM64_INSTR_PT(528)
     OR ROM64_INSTR_PT(529) OR ROM64_INSTR_PT(537)
     OR ROM64_INSTR_PT(542) OR ROM64_INSTR_PT(550)
     OR ROM64_INSTR_PT(560) OR ROM64_INSTR_PT(566)
     OR ROM64_INSTR_PT(573) OR ROM64_INSTR_PT(581)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(607)
     OR ROM64_INSTR_PT(621) OR ROM64_INSTR_PT(661)
     OR ROM64_INSTR_PT(698) OR ROM64_INSTR_PT(706)
     OR ROM64_INSTR_PT(790) OR ROM64_INSTR_PT(823)
     OR ROM64_INSTR_PT(854));
MQQ936:SEL6_10(1) <= 
    (ROM64_INSTR_PT(1) OR ROM64_INSTR_PT(3)
     OR ROM64_INSTR_PT(40) OR ROM64_INSTR_PT(54)
     OR ROM64_INSTR_PT(67) OR ROM64_INSTR_PT(69)
     OR ROM64_INSTR_PT(78) OR ROM64_INSTR_PT(82)
     OR ROM64_INSTR_PT(95) OR ROM64_INSTR_PT(107)
     OR ROM64_INSTR_PT(120) OR ROM64_INSTR_PT(182)
     OR ROM64_INSTR_PT(188) OR ROM64_INSTR_PT(256)
     OR ROM64_INSTR_PT(267) OR ROM64_INSTR_PT(287)
     OR ROM64_INSTR_PT(336) OR ROM64_INSTR_PT(346)
     OR ROM64_INSTR_PT(350) OR ROM64_INSTR_PT(354)
     OR ROM64_INSTR_PT(358) OR ROM64_INSTR_PT(380)
     OR ROM64_INSTR_PT(407) OR ROM64_INSTR_PT(431)
     OR ROM64_INSTR_PT(436) OR ROM64_INSTR_PT(459)
     OR ROM64_INSTR_PT(463) OR ROM64_INSTR_PT(487)
     OR ROM64_INSTR_PT(529) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(540) OR ROM64_INSTR_PT(580)
     OR ROM64_INSTR_PT(605) OR ROM64_INSTR_PT(640)
     OR ROM64_INSTR_PT(652) OR ROM64_INSTR_PT(658)
     OR ROM64_INSTR_PT(694) OR ROM64_INSTR_PT(697)
     OR ROM64_INSTR_PT(708) OR ROM64_INSTR_PT(715)
     OR ROM64_INSTR_PT(718) OR ROM64_INSTR_PT(720)
     OR ROM64_INSTR_PT(726) OR ROM64_INSTR_PT(727)
     OR ROM64_INSTR_PT(740) OR ROM64_INSTR_PT(769)
     OR ROM64_INSTR_PT(857) OR ROM64_INSTR_PT(864)
    );
MQQ937:SEL11_15(0) <= 
    (ROM64_INSTR_PT(37) OR ROM64_INSTR_PT(135)
     OR ROM64_INSTR_PT(193) OR ROM64_INSTR_PT(232)
     OR ROM64_INSTR_PT(248) OR ROM64_INSTR_PT(291)
     OR ROM64_INSTR_PT(373) OR ROM64_INSTR_PT(384)
     OR ROM64_INSTR_PT(438) OR ROM64_INSTR_PT(447)
     OR ROM64_INSTR_PT(465) OR ROM64_INSTR_PT(593)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(741)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(829)
    );
MQQ938:SEL11_15(1) <= 
    (ROM64_INSTR_PT(24) OR ROM64_INSTR_PT(27)
     OR ROM64_INSTR_PT(37) OR ROM64_INSTR_PT(44)
     OR ROM64_INSTR_PT(48) OR ROM64_INSTR_PT(59)
     OR ROM64_INSTR_PT(62) OR ROM64_INSTR_PT(63)
     OR ROM64_INSTR_PT(85) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(105) OR ROM64_INSTR_PT(115)
     OR ROM64_INSTR_PT(123) OR ROM64_INSTR_PT(130)
     OR ROM64_INSTR_PT(133) OR ROM64_INSTR_PT(140)
     OR ROM64_INSTR_PT(141) OR ROM64_INSTR_PT(151)
     OR ROM64_INSTR_PT(164) OR ROM64_INSTR_PT(189)
     OR ROM64_INSTR_PT(192) OR ROM64_INSTR_PT(193)
     OR ROM64_INSTR_PT(200) OR ROM64_INSTR_PT(220)
     OR ROM64_INSTR_PT(232) OR ROM64_INSTR_PT(234)
     OR ROM64_INSTR_PT(250) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(266) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(291) OR ROM64_INSTR_PT(303)
     OR ROM64_INSTR_PT(323) OR ROM64_INSTR_PT(354)
     OR ROM64_INSTR_PT(356) OR ROM64_INSTR_PT(373)
     OR ROM64_INSTR_PT(386) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(418) OR ROM64_INSTR_PT(423)
     OR ROM64_INSTR_PT(432) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(444)
     OR ROM64_INSTR_PT(452) OR ROM64_INSTR_PT(465)
     OR ROM64_INSTR_PT(492) OR ROM64_INSTR_PT(516)
     OR ROM64_INSTR_PT(524) OR ROM64_INSTR_PT(528)
     OR ROM64_INSTR_PT(547) OR ROM64_INSTR_PT(550)
     OR ROM64_INSTR_PT(560) OR ROM64_INSTR_PT(573)
     OR ROM64_INSTR_PT(577) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(593) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(607) OR ROM64_INSTR_PT(621)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(634)
     OR ROM64_INSTR_PT(665) OR ROM64_INSTR_PT(698)
     OR ROM64_INSTR_PT(706) OR ROM64_INSTR_PT(717)
     OR ROM64_INSTR_PT(718) OR ROM64_INSTR_PT(734)
     OR ROM64_INSTR_PT(790) OR ROM64_INSTR_PT(806)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(824)
     OR ROM64_INSTR_PT(828) OR ROM64_INSTR_PT(840)
     OR ROM64_INSTR_PT(844) OR ROM64_INSTR_PT(849)
    );
MQQ939:SEL16_20(0) <= 
    (ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(135)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(258)
     OR ROM64_INSTR_PT(260) OR ROM64_INSTR_PT(355)
     OR ROM64_INSTR_PT(447) OR ROM64_INSTR_PT(533)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(829)
    );
MQQ940:SEL16_20(1) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(12)
     OR ROM64_INSTR_PT(16) OR ROM64_INSTR_PT(40)
     OR ROM64_INSTR_PT(46) OR ROM64_INSTR_PT(48)
     OR ROM64_INSTR_PT(69) OR ROM64_INSTR_PT(74)
     OR ROM64_INSTR_PT(82) OR ROM64_INSTR_PT(87)
     OR ROM64_INSTR_PT(95) OR ROM64_INSTR_PT(100)
     OR ROM64_INSTR_PT(107) OR ROM64_INSTR_PT(126)
     OR ROM64_INSTR_PT(133) OR ROM64_INSTR_PT(135)
     OR ROM64_INSTR_PT(137) OR ROM64_INSTR_PT(141)
     OR ROM64_INSTR_PT(159) OR ROM64_INSTR_PT(164)
     OR ROM64_INSTR_PT(200) OR ROM64_INSTR_PT(204)
     OR ROM64_INSTR_PT(225) OR ROM64_INSTR_PT(251)
     OR ROM64_INSTR_PT(266) OR ROM64_INSTR_PT(267)
     OR ROM64_INSTR_PT(279) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(300) OR ROM64_INSTR_PT(319)
     OR ROM64_INSTR_PT(321) OR ROM64_INSTR_PT(336)
     OR ROM64_INSTR_PT(354) OR ROM64_INSTR_PT(355)
     OR ROM64_INSTR_PT(362) OR ROM64_INSTR_PT(379)
     OR ROM64_INSTR_PT(398) OR ROM64_INSTR_PT(413)
     OR ROM64_INSTR_PT(423) OR ROM64_INSTR_PT(444)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(447)
     OR ROM64_INSTR_PT(452) OR ROM64_INSTR_PT(470)
     OR ROM64_INSTR_PT(496) OR ROM64_INSTR_PT(513)
     OR ROM64_INSTR_PT(524) OR ROM64_INSTR_PT(528)
     OR ROM64_INSTR_PT(529) OR ROM64_INSTR_PT(541)
     OR ROM64_INSTR_PT(550) OR ROM64_INSTR_PT(560)
     OR ROM64_INSTR_PT(561) OR ROM64_INSTR_PT(566)
     OR ROM64_INSTR_PT(572) OR ROM64_INSTR_PT(573)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(607)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(621)
     OR ROM64_INSTR_PT(634) OR ROM64_INSTR_PT(648)
     OR ROM64_INSTR_PT(661) OR ROM64_INSTR_PT(698)
     OR ROM64_INSTR_PT(706) OR ROM64_INSTR_PT(717)
     OR ROM64_INSTR_PT(729) OR ROM64_INSTR_PT(773)
     OR ROM64_INSTR_PT(790) OR ROM64_INSTR_PT(798)
     OR ROM64_INSTR_PT(829) OR ROM64_INSTR_PT(838)
    );
MQQ941:SEL21_25(0) <= 
    (ROM64_INSTR_PT(197));
MQQ942:SEL21_25(1) <= 
    (ROM64_INSTR_PT(16) OR ROM64_INSTR_PT(46)
     OR ROM64_INSTR_PT(48) OR ROM64_INSTR_PT(63)
     OR ROM64_INSTR_PT(74) OR ROM64_INSTR_PT(87)
     OR ROM64_INSTR_PT(141) OR ROM64_INSTR_PT(200)
     OR ROM64_INSTR_PT(225) OR ROM64_INSTR_PT(266)
     OR ROM64_INSTR_PT(321) OR ROM64_INSTR_PT(354)
     OR ROM64_INSTR_PT(362) OR ROM64_INSTR_PT(423)
     OR ROM64_INSTR_PT(452) OR ROM64_INSTR_PT(470)
     OR ROM64_INSTR_PT(515) OR ROM64_INSTR_PT(528)
     OR ROM64_INSTR_PT(541) OR ROM64_INSTR_PT(550)
     OR ROM64_INSTR_PT(560) OR ROM64_INSTR_PT(572)
     OR ROM64_INSTR_PT(573) OR ROM64_INSTR_PT(634)
     OR ROM64_INSTR_PT(652) OR ROM64_INSTR_PT(706)
     OR ROM64_INSTR_PT(718) OR ROM64_INSTR_PT(729)
     OR ROM64_INSTR_PT(734) OR ROM64_INSTR_PT(790)
    );
MQQ943:SEL26_30 <= 
    (ROM64_INSTR_PT(16) OR ROM64_INSTR_PT(46)
     OR ROM64_INSTR_PT(48) OR ROM64_INSTR_PT(63)
     OR ROM64_INSTR_PT(74) OR ROM64_INSTR_PT(87)
     OR ROM64_INSTR_PT(141) OR ROM64_INSTR_PT(200)
     OR ROM64_INSTR_PT(225) OR ROM64_INSTR_PT(266)
     OR ROM64_INSTR_PT(321) OR ROM64_INSTR_PT(354)
     OR ROM64_INSTR_PT(362) OR ROM64_INSTR_PT(423)
     OR ROM64_INSTR_PT(452) OR ROM64_INSTR_PT(470)
     OR ROM64_INSTR_PT(515) OR ROM64_INSTR_PT(528)
     OR ROM64_INSTR_PT(541) OR ROM64_INSTR_PT(550)
     OR ROM64_INSTR_PT(560) OR ROM64_INSTR_PT(572)
     OR ROM64_INSTR_PT(573) OR ROM64_INSTR_PT(634)
     OR ROM64_INSTR_PT(652) OR ROM64_INSTR_PT(706)
     OR ROM64_INSTR_PT(718) OR ROM64_INSTR_PT(729)
     OR ROM64_INSTR_PT(734) OR ROM64_INSTR_PT(790)
    );
MQQ944:SEL31 <= 
    (ROM64_INSTR_PT(16) OR ROM64_INSTR_PT(46)
     OR ROM64_INSTR_PT(63) OR ROM64_INSTR_PT(74)
     OR ROM64_INSTR_PT(87) OR ROM64_INSTR_PT(141)
     OR ROM64_INSTR_PT(200) OR ROM64_INSTR_PT(266)
     OR ROM64_INSTR_PT(321) OR ROM64_INSTR_PT(350)
     OR ROM64_INSTR_PT(354) OR ROM64_INSTR_PT(358)
     OR ROM64_INSTR_PT(362) OR ROM64_INSTR_PT(423)
     OR ROM64_INSTR_PT(452) OR ROM64_INSTR_PT(470)
     OR ROM64_INSTR_PT(541) OR ROM64_INSTR_PT(542)
     OR ROM64_INSTR_PT(560) OR ROM64_INSTR_PT(561)
     OR ROM64_INSTR_PT(573) OR ROM64_INSTR_PT(634)
     OR ROM64_INSTR_PT(652) OR ROM64_INSTR_PT(697)
     OR ROM64_INSTR_PT(706) OR ROM64_INSTR_PT(715)
     OR ROM64_INSTR_PT(718) OR ROM64_INSTR_PT(729)
     OR ROM64_INSTR_PT(790) OR ROM64_INSTR_PT(823)
    );
MQQ945:CR_BF2FXM <= 
    (ROM64_INSTR_PT(717));
MQQ946:SKIP_COND <= 
    (ROM64_INSTR_PT(23) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(81) OR ROM64_INSTR_PT(88)
     OR ROM64_INSTR_PT(91) OR ROM64_INSTR_PT(127)
     OR ROM64_INSTR_PT(298) OR ROM64_INSTR_PT(330)
     OR ROM64_INSTR_PT(331) OR ROM64_INSTR_PT(335)
     OR ROM64_INSTR_PT(344) OR ROM64_INSTR_PT(369)
     OR ROM64_INSTR_PT(489) OR ROM64_INSTR_PT(662)
     OR ROM64_INSTR_PT(667) OR ROM64_INSTR_PT(677)
     OR ROM64_INSTR_PT(684) OR ROM64_INSTR_PT(725)
     OR ROM64_INSTR_PT(744) OR ROM64_INSTR_PT(745)
     OR ROM64_INSTR_PT(746) OR ROM64_INSTR_PT(747)
     OR ROM64_INSTR_PT(748) OR ROM64_INSTR_PT(750)
     OR ROM64_INSTR_PT(754) OR ROM64_INSTR_PT(755)
     OR ROM64_INSTR_PT(756) OR ROM64_INSTR_PT(765)
     OR ROM64_INSTR_PT(776) OR ROM64_INSTR_PT(782)
     OR ROM64_INSTR_PT(783) OR ROM64_INSTR_PT(784)
     OR ROM64_INSTR_PT(792) OR ROM64_INSTR_PT(795)
     OR ROM64_INSTR_PT(796) OR ROM64_INSTR_PT(804)
     OR ROM64_INSTR_PT(817) OR ROM64_INSTR_PT(819)
     OR ROM64_INSTR_PT(820) OR ROM64_INSTR_PT(821)
     OR ROM64_INSTR_PT(827) OR ROM64_INSTR_PT(842)
     OR ROM64_INSTR_PT(859) OR ROM64_INSTR_PT(867)
    );
MQQ947:SKIP_ZERO <= 
    (ROM64_INSTR_PT(301) OR ROM64_INSTR_PT(319)
     OR ROM64_INSTR_PT(393) OR ROM64_INSTR_PT(436)
     OR ROM64_INSTR_PT(487) OR ROM64_INSTR_PT(496)
     OR ROM64_INSTR_PT(778));
MQQ948:LOOP_ADDR(0) <= 
    (ROM64_INSTR_PT(235) OR ROM64_INSTR_PT(289)
     OR ROM64_INSTR_PT(301) OR ROM64_INSTR_PT(317)
     OR ROM64_INSTR_PT(328) OR ROM64_INSTR_PT(373)
     OR ROM64_INSTR_PT(479) OR ROM64_INSTR_PT(526)
     OR ROM64_INSTR_PT(674) OR ROM64_INSTR_PT(692)
     OR ROM64_INSTR_PT(700) OR ROM64_INSTR_PT(732)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(777)
     OR ROM64_INSTR_PT(778) OR ROM64_INSTR_PT(784)
     OR ROM64_INSTR_PT(837) OR ROM64_INSTR_PT(861)
     OR ROM64_INSTR_PT(866) OR ROM64_INSTR_PT(867)
    );
MQQ949:LOOP_ADDR(1) <= 
    (ROM64_INSTR_PT(289) OR ROM64_INSTR_PT(479)
     OR ROM64_INSTR_PT(526) OR ROM64_INSTR_PT(674)
     OR ROM64_INSTR_PT(732) OR ROM64_INSTR_PT(777)
     OR ROM64_INSTR_PT(784) OR ROM64_INSTR_PT(833)
     OR ROM64_INSTR_PT(837) OR ROM64_INSTR_PT(859)
     OR ROM64_INSTR_PT(867));
MQQ950:LOOP_ADDR(2) <= 
    (ROM64_INSTR_PT(393) OR ROM64_INSTR_PT(449)
     OR ROM64_INSTR_PT(486) OR ROM64_INSTR_PT(700)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(748)
     OR ROM64_INSTR_PT(754) OR ROM64_INSTR_PT(764)
    );
MQQ951:LOOP_ADDR(3) <= 
    (ROM64_INSTR_PT(317) OR ROM64_INSTR_PT(328)
     OR ROM64_INSTR_PT(501) OR ROM64_INSTR_PT(672)
     OR ROM64_INSTR_PT(688) OR ROM64_INSTR_PT(700)
     OR ROM64_INSTR_PT(707) OR ROM64_INSTR_PT(725)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(765)
     OR ROM64_INSTR_PT(767) OR ROM64_INSTR_PT(777)
     OR ROM64_INSTR_PT(836) OR ROM64_INSTR_PT(837)
     OR ROM64_INSTR_PT(859) OR ROM64_INSTR_PT(867)
     OR ROM64_INSTR_PT(878));
MQQ952:LOOP_ADDR(4) <= 
    (ROM64_INSTR_PT(37) OR ROM64_INSTR_PT(289)
     OR ROM64_INSTR_PT(301) OR ROM64_INSTR_PT(328)
     OR ROM64_INSTR_PT(373) OR ROM64_INSTR_PT(400)
     OR ROM64_INSTR_PT(421) OR ROM64_INSTR_PT(449)
     OR ROM64_INSTR_PT(479) OR ROM64_INSTR_PT(700)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(748)
     OR ROM64_INSTR_PT(750) OR ROM64_INSTR_PT(754)
     OR ROM64_INSTR_PT(762) OR ROM64_INSTR_PT(784)
     OR ROM64_INSTR_PT(837) OR ROM64_INSTR_PT(866)
     OR ROM64_INSTR_PT(867));
MQQ953:LOOP_ADDR(5) <= 
    (ROM64_INSTR_PT(37) OR ROM64_INSTR_PT(235)
     OR ROM64_INSTR_PT(289) OR ROM64_INSTR_PT(421)
     OR ROM64_INSTR_PT(449) OR ROM64_INSTR_PT(526)
     OR ROM64_INSTR_PT(688) OR ROM64_INSTR_PT(725)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(764)
     OR ROM64_INSTR_PT(772) OR ROM64_INSTR_PT(861)
     OR ROM64_INSTR_PT(866));
MQQ954:LOOP_ADDR(6) <= 
    (ROM64_INSTR_PT(37) OR ROM64_INSTR_PT(163)
     OR ROM64_INSTR_PT(289) OR ROM64_INSTR_PT(317)
     OR ROM64_INSTR_PT(373) OR ROM64_INSTR_PT(486)
     OR ROM64_INSTR_PT(672) OR ROM64_INSTR_PT(696)
     OR ROM64_INSTR_PT(700) OR ROM64_INSTR_PT(748)
     OR ROM64_INSTR_PT(750) OR ROM64_INSTR_PT(764)
     OR ROM64_INSTR_PT(767) OR ROM64_INSTR_PT(833)
     OR ROM64_INSTR_PT(837) OR ROM64_INSTR_PT(859)
     OR ROM64_INSTR_PT(861) OR ROM64_INSTR_PT(868)
    );
MQQ955:LOOP_ADDR(7) <= 
    (ROM64_INSTR_PT(37) OR ROM64_INSTR_PT(289)
     OR ROM64_INSTR_PT(301) OR ROM64_INSTR_PT(317)
     OR ROM64_INSTR_PT(328) OR ROM64_INSTR_PT(400)
     OR ROM64_INSTR_PT(421) OR ROM64_INSTR_PT(486)
     OR ROM64_INSTR_PT(651) OR ROM64_INSTR_PT(672)
     OR ROM64_INSTR_PT(674) OR ROM64_INSTR_PT(692)
     OR ROM64_INSTR_PT(725) OR ROM64_INSTR_PT(732)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(748)
     OR ROM64_INSTR_PT(777) OR ROM64_INSTR_PT(861)
     OR ROM64_INSTR_PT(867));
MQQ956:LOOP_ADDR(8) <= 
    (ROM64_INSTR_PT(400) OR ROM64_INSTR_PT(421)
     OR ROM64_INSTR_PT(449) OR ROM64_INSTR_PT(479)
     OR ROM64_INSTR_PT(486) OR ROM64_INSTR_PT(672)
     OR ROM64_INSTR_PT(696) OR ROM64_INSTR_PT(700)
     OR ROM64_INSTR_PT(707) OR ROM64_INSTR_PT(725)
     OR ROM64_INSTR_PT(748) OR ROM64_INSTR_PT(750)
     OR ROM64_INSTR_PT(754) OR ROM64_INSTR_PT(762)
     OR ROM64_INSTR_PT(764) OR ROM64_INSTR_PT(777)
     OR ROM64_INSTR_PT(861) OR ROM64_INSTR_PT(866)
    );
MQQ957:LOOP_ADDR(9) <= 
    (ROM64_INSTR_PT(301) OR ROM64_INSTR_PT(317)
     OR ROM64_INSTR_PT(328) OR ROM64_INSTR_PT(373)
     OR ROM64_INSTR_PT(393) OR ROM64_INSTR_PT(449)
     OR ROM64_INSTR_PT(486) OR ROM64_INSTR_PT(692)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(764)
     OR ROM64_INSTR_PT(772) OR ROM64_INSTR_PT(778)
     OR ROM64_INSTR_PT(784) OR ROM64_INSTR_PT(836)
     OR ROM64_INSTR_PT(837) OR ROM64_INSTR_PT(861)
    );
MQQ958:LOOP_INIT(0) <= 
    (ROM64_INSTR_PT(235) OR ROM64_INSTR_PT(369)
     OR ROM64_INSTR_PT(398) OR ROM64_INSTR_PT(572)
     OR ROM64_INSTR_PT(673) OR ROM64_INSTR_PT(692)
     OR ROM64_INSTR_PT(783) OR ROM64_INSTR_PT(795)
     OR ROM64_INSTR_PT(810) OR ROM64_INSTR_PT(817)
     OR ROM64_INSTR_PT(821) OR ROM64_INSTR_PT(837)
     OR ROM64_INSTR_PT(859) OR ROM64_INSTR_PT(867)
    );
MQQ959:LOOP_INIT(1) <= 
    (ROM64_INSTR_PT(890));
MQQ960:LOOP_INIT(2) <= 
    (ROM64_INSTR_PT(783) OR ROM64_INSTR_PT(817)
     OR ROM64_INSTR_PT(859) OR ROM64_INSTR_PT(867)
    );
MQQ961:EP <= 
    (ROM64_INSTR_PT(44) OR ROM64_INSTR_PT(59)
     OR ROM64_INSTR_PT(115) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(279) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(356) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(398) OR ROM64_INSTR_PT(432)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(524) OR ROM64_INSTR_PT(561)
    );

end generate;
--32-bit core
c32: if (regmode = 5) generate
begin

ROM64_INSTR_PT  <=  (others => '0');
rom_unused  <=  or_reduce(ROM64_INSTR_PT);
--
-- Final Table Listing
--      *INPUTS*========*OUTPUTS*===============================================================================================*
--      |               |                                                                                                       |
--      | rom_addr_l2   | template                         ucode_end                                                            |
--      | |             | |                                | ucode_end_early                                                    |
--      | |             | |                                | | loop_begin                                                       |
--      | |             | |                                | | | loop_end                                                       |
--      | |             | |                                | | | | count_src                                                    | -- Can DC if not (loop_begin or loop_end)
--      | |             | |                                | | | | |                                                            |
--      | |             | |                                | | | | |    extRT                                                   |
--      | |             | |                                | | | | |    | extS1                                                 |
--      | |             | |                                | | | | |    | | extS2                                               |
--      | |             | |                                | | | | |    | | | extS3                                             |
--      | |             | |                                | | | | |    | | | |                                                 |
--      | |             | |                                | | | | |    | | | |  sel0_5                                         |
--      | |             | |                                | | | | |    | | | |  | sel6_10                                      |
--      | |             | |                                | | | | |    | | | |  | |  sel11_15                                  |
--      | |             | |                                | | | | |    | | | |  | |  |  sel16_20                               |
--      | |             | |                                | | | | |    | | | |  | |  |  |  sel21_25                            |
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  sel26_30                         |
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | sel31                          |
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | |                              |
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | |  cr_bf2fxm                   |
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | skip_cond                 |
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | skip_zero               | -- Can DC if loop_begin not set
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | | loop_addr             | -- Can DC if loop_end not set
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | | |          loop_init  | -- 1 less than # of times to loop; Can DC if not loop_end or not count_src=111
--      | |             | |                                | | | | |    | | | |  | |  |  |  |  | |  | | | |          |   ep     |
--      | |             | |         1111111111222222222233 | | | | |    | | | |  | |  |  |  |  | |  | | | |          |   |      |
--      | 0123456789    | 01234567890123456789012345678901 | | | | 012  | | | |  | 01 01 01 01 | |  | | | 0123456789 012 |      |
--      *TYPE*==========+=======================================================================================================+
--      | PPPPPPPPPP    | SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSS S S S S SSS  S S S S  S SS SS SS SS S S  S S S SSSSSSSSSS SSS S      |
--      *POLARITY*----->| ++++++++++++++++++++++++++++++++ + + + + +++  + + + +  + ++ ++ ++ ++ + +  + + + ++++++++++ +++ +      |
--      *PHASE*-------->| TTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTT T T T T TTT  T T T T  T TT TT TT TT T T  T T T TTTTTTTTTT TTT T      |
--      *OPTIMIZE*----->|  AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA B B B B CCC  X X X X  X XX XX XX XX X X  X X X XXXXXXXXXX XYX X       |
--      *TERMS*=========+=======================================================================================================+
--    1 | -100000000    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--    2 | 0-11000000    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--    3 | 10-1000000    | .1...1....1.............1.1.111. . . . . ...  1 1 . .  . .. .. .1 .. . .  . . . .......... ... .      |
--    4 | 000-000000    | ..111...........111111111111111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--    5 | 110-000000    | .11111....1..........1.1111111.. . . . . ...  . . . .  . .. .. 1. .. . .  . . . .......... ... .      |
--    6 | 011-000000    | .11111...11...1...........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--    7 | -0-0100000    | .11111................1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--    8 | 0001100000    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--    9 | 01-1100000    | .1.1.1..........1....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   10 | -01-100000    | .1.1.1...1....1......11.1.11.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   11 | -000-00000    | ................................ . . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   12 | 11-0-00000    | .....1...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   13 | 0001010000    | .11111....1.............1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   14 | 0-11010000    | .11111...11...11...1..1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   15 | 10-1010000    | ................................ . . . . ...  . . . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   16 | 0-00110000    | .1.1......1...1.11..........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   17 | -1-0110000    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   18 | 0-11110000    | ..111.....1.....1111............ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   19 | 10--110000    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . 1..11..1.1 ... .      |
--   20 | 01--110000    | .1.1.1........1.1111111..111..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   21 | 0000-10000    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   22 | 1101-10000    | ................................ . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   23 | 011--10000    | .1111....1....1....1.111.11..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   24 | 11-00-0000    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   25 | 00010-0000    | ................................ . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   26 | 01001-0000    | .1.1.1........111111....1.11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   27 | 10-01-0000    | ..111........................1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   28 | 11011-0000    | 1..11....1...................... . . . . ...  . 1 . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   29 | 011-1-0000    | ..1.1.................1.1.1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   30 | 1-1-1-0000    | .............................1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   31 | 1001--0000    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   32 | 101---0000    | .1.1......1...1.11..........1.1. . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   33 | 111---0000    | 1..111..............1.....11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   34 | 0-00001000    | ..............111111....1....... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   35 | --10001000    | .1111....1....1.....1111111..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   36 | 10-1001000    | ................................ . . . . ...  . 1 1 .  . .. 11 .. .. . .  . . . 1...1111.1 ... .      |
--   37 | 110-001000    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   38 | -01-001000    | ..111.....1.....11111111........ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   39 | -100101000    | .11111.............1......111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   40 | 11-0101000    | ................................ . . . . ...  1 . . .  . 11 .. .1 .. . .  . . . .......... ... .      |
--   41 | 0001101000    | .11111....1.............1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   42 | 0-11101000    | .11111...11...1....11....1.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   43 | 01-1101000    | .1111............1...11...1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   44 | 000-101000    | ................................ . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... 1      |
--   45 | 111-101000    | 1..111...11........11...1.111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   46 | 0000-01000    | ................................ . . . . ...  . . . .  . .. .. .1 .1 1 .  . . . .......... ... .      |
--   47 | -11--01000    | ................................ . . . . ...  1 1 1 1  . .. .. .. .. . .  . . . .......... ... .      |
--   48 | 0001011000    | ................................ . . . . ...  . . . .  . .. .1 .1 .1 1 .  . . . .......... ... .      |
--   49 | 0-11011000    | .1.1.1..........11111.....11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   50 | 01-1011000    | .1........................1...1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   51 | 00-0111000    | .1...1....1.............1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   52 | 110-111000    | .1.1.1....1...1...........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   53 | 0-1-111000    | .11111...11...11...1..1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   54 | 0100-11000    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   55 | 1101-11000    | .1.......1....1.11............1. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   56 | 101--11000    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   57 | 011--11000    | .11111....1....1...1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   58 | --1--11000    | ................................ . . . . ...  . 1 . 1  . .. .. .. .. . .  . . . 1.1111.1.1 ... .      |
--   59 | 01000-1000    | .1.1.1....................11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   60 | -0100-1000    | .........1...........1....1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   61 | 00001-1000    | ................................ . . . . ...  . . . .  . .. .1 .. .. . 1  . . . .......... ... 1      |
--   62 | 00-01-1000    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   63 | 10011-1000    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   64 | 11011-1000    | ................................ . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   65 | 000000-000    | ................................ . . . . ...  . . . .  . .. .1 .. .1 1 1  . . . .......... ... .      |
--   66 | -10000-000    | .1.1.1....................11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   67 | -01000-000    | .1.1.1........1.1...........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   68 | 10-000-000    | 1...1........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   69 | 10-010-000    | ................................ . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   70 | 1--010-000    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   71 | 01-110-000    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   72 | 101--0-000    | .11111....................111... . . . . ...  1 . . .  . 11 .. .1 .. . .  . . . .......... ... .      |
--   73 | 000001-000    | .1.1.1...1....1..1...1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   74 | 0-1011-000    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   75 | -------000    | ................................ . . . . 1..  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   76 | 0001000100    | 1...1.....1..................... . . . . ...  . . . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   77 | 1101000100    | .1.1......1...1.1...........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   78 | 0-11000100    | ...1.................11...1..11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   79 | 01-1000100    | .1111.........111111....1.....1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   80 | 011-000100    | .1111............1...11...1...1. . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   81 | 10--000100    | ..1.1..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   82 | 11-0100100    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   83 | 0001100100    | .11111....................111... . . . . ...  . . . .  . 11 .. .1 .. . .  . . . .......... ... .      |
--   84 | 0-11100100    | .1.1.1.........11....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   85 | 1-1-100100    | 1..111...11...1....1......111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   86 | 10--100100    | ................................ . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   87 | 0000-00100    | .1.1.1...1....1..1...1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   88 | 10-0-00100    | ................................ . . . . ...  . . . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   89 | 1101-00100    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   90 | 11-0010100    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   91 | 0001010100    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   92 | 010-010100    | .1111.........11..........1...1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   93 | -01-010100    | .1.1.1...1....1......1111.1111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   94 | 0-00110100    | ................................ . . . . ...  1 . . .  . 11 .. .1 .. . .  . . . .......... ... .      |
--   95 | -1-0110100    | ..111.....1.....1111111111111..1 . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   96 | 000-110100    | .1...1....................11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   97 | 01--110100    | .1111....1....1...11.11..11..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   98 | 0-00-10100    | ..111.......................1... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   99 | 0001-10100    | .1.1......1...1.11..........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   100 | 1101-10100    | .1...1...1.............11.1.111. . . . . ...  . 1 . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   101 | 011--10100    | .11111.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   102 | 01000-0100    | .11111...1.....1...11.....111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   103 | -0100-0100    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   104 | 10-01-0100    | ...............................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   105 | 11011-0100    | .1111....1....1.11............1. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   106 | 101---0100    | .1...1...1..............1.1.111. . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   107 | 111---0100    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   108 | 0001001100    | ................................ . . . . ...  1 . . .  . 11 .. .1 .. . .  . . . .......... ... .      |
--   109 | -001001100    | .11111....................111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   110 | --11001100    | .11111.............1......11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   111 | 01-1001100    | .1111.........111.1....1......1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   112 | -1-1001100    | .................1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   113 | 00-0101100    | 1...1.....1..................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   114 | 10-0101100    | .1.1......1...1.1.....1....1111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   115 | 01-0101100    | .1.1.1........111....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   116 | 11-0101100    | ...1.1..................1.1.111. . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... 1      |
--   117 | 01-1101100    | .11111...11....1..........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   118 | 0-1-101100    | .1.1.1....1...1.1....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   119 | 011--01100    | .1.1.1........1.1111111..111..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   120 | 11-0011100    | 1...1....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   121 | --11011100    | ................................ . . . . ...  1 . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   122 | 01-1011100    | .1111..........111....1.......1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   123 | -1-1111100    | ..........1....1................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   124 | 110-111100    | .11111...1.............11.1.111. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   125 | 0-1-111100    | ..........1...1..........1..1... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   126 | 11--111100    | ................................ . . . . ...  . . . 1  . .. .. .1 .. . .  . . . .......... ... .      |
--   127 | 0000-11100    | .1.1......1...1.11..........111. . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   128 | 0001-11100    | 1...1.....1..................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   129 | 11-1-11100    | ................................ . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   130 | 011--11100    | .11111...11...1...........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   131 | 10-00-1100    | ...1.1................1....1.1.. . . . . ...  1 . . .  . .. .1 .1 .. . .  . . . .......... ... .      |
--   132 | -1110-1100    | 1........................1..11.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   133 | 1-1-0-1100    | ................................ . . . . ...  1 . . 1  . .. 1. 11 .. . .  . . . .......... ... .      |
--   134 | 00011-1100    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   135 | 1-011-1100    | .1...1...1.............11.1.111. . . . . ...  . 1 . 1  . .. .. .1 .. . .  . . . .......... ... 1      |
--   136 | 0---1-1100    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . ...11.1.1. ... .      |
--   137 | -01-00-100    | ................................ . . . . ...  . 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   138 | 11-010-100    | ....1.....1...1................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   139 | 101--0-100    | .11111....1.............1.1.111. . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   140 | 000001-100    | ................................ . . . . ...  . . . .  . .. .1 .1 .1 1 1  . . . .......... ... .      |
--   141 | 010001-100    | .11111...1.....1...11.....111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   142 | 1-1-01-100    | 1...11...11.............11111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   143 | 01-011-100    | .....1....1...1....1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   144 | 0-1111-100    | .11111.............1......11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   145 | -010-1-100    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   146 | 10-0-1-100    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   147 | 11-0000-00    | ..111..........................1 . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   148 | -010100-00    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   149 | ---0100-00    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   150 | -010010-00    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   151 | 10--010-00    | ..111........................... . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   152 | --1---0-00    | ................................ . . . . ...  1 . 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   153 | 0000001-00    | .11111....1.............1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   154 | -010001-00    | .........1...........1....1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   155 | 10-1001-00    | ...111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   156 | ----001-00    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   157 | 0-1--01-00    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   158 | 01-1111-00    | .11111.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   159 | 11-1111-00    | 1...11.........1........111111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   160 | 100-111-00    | ................................ . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   161 | -11-111-00    | ................................ . . . . ...  1 . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   162 | 1001-11-00    | 1..11....1.....................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   163 | 011-1-1-00    | .11111.........1....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   164 | 10-001--00    | .1.1.1................1....1.1.. . . . . ...  1 . . .  . .. .1 .1 .. . .  . . . .......... ... .      |
--   165 | 01-011--00    | .1111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   166 | 1101-1--00    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   167 | 0-1-1---00    | ................................ . . . . ...  . 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   168 | -101----00    | ................................ . . . . ...  1 . . 1  . .. .. .. .. . .  . . . .......... 1.1 .      |
--   169 | 1101000010    | .1.1.1....1...1...........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   170 | 0-11000010    | .1...1.........1........11.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   171 | 10-1000010    | .1.1......1...1.1.....1....1111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   172 | 011-000010    | .1111....1....1...1..11.111..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   173 | 11-0100010    | ...11.....1....1.1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   174 | 0-11100010    | ..111....11...11..........1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   175 | 0000-00010    | 1...1....1.....................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   176 | 1-1--00010    | 1..111...1................11..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   177 | -010010010    | 1..11....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   178 | -1-0110010    | ...11..............1.1...1.1.... . . . . ...  . . 1 .  . .1 .. .. .. . .  . . . .......... ... .      |
--   179 | 00-1110010    | .1.1.1...1....1......111.1111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   180 | -11-110010    | 1..111...11...............11..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   181 | 01--110010    | ...111...11...1...........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   182 | -110-10010    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   183 | 11-0-10010    | .1...1....1.............1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   184 | 0001-10010    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   185 | 1101-10010    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   186 | 011--10010    | .1111...........11...11...1...1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   187 | 01000-0010    | ..1111...1....1..1.1.1.1.1.1.1.1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   188 | 11-00-0010    | ................................ . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   189 | 0-110-0010    | ..111.....1.....11.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   190 | 1-1-0-0010    | ................................ . . . . ...  1 . . 1  . .. .1 .. .. . .  . . . .......... ... .      |
--   191 | -0--0-0010    | ................................ . . . . ...  . . 1 .  . .. .. .. .. . .  . . . .........1 ... .      |
--   192 | 01001-0010    | .11111...1................111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   193 | 00011-0010    | .11.1....1...................... . . . . ...  . 1 . .  . .. 11 .. .. . .  . . . .......... ... .      |
--   194 | 11011-0010    | ...111....1..........1.11111111. . . . . ...  . . . .  . .. .. 1. .. . .  . . . .......... ... .      |
--   195 | 1--11-0010    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   196 | 011-1-0010    | .1...1........1.....1.1..1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   197 | 111-1-0010    | ................................ . . . . ...  1 1 . .  . .. .. .. 1. . .  . . . .......... ... .      |
--   198 | 101---0010    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   199 | 0-00001010    | .11111...1................111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   200 | 1--0001010    | .1.1......1...1.11..........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   201 | 1101001010    | ................................ 1 . . . ...  . . . .  . 1. .1 .1 .1 1 1  . . . .......... ... .      |
--   202 | 00-1001010    | .1.1.1...1....1......111..111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   203 | 011-001010    | .11111....1....1...1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   204 | 10--001010    | .....1....1.............1.1.111. . . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   205 | 0100101010    | .11111.............11.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   206 | 0-11101010    | .11111.............1.1....11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   207 | 01-1101010    | .11111.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   208 | 110-101010    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   209 | 0001-01010    | .1111....1....1.11............1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   210 | 1-01-01010    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   211 | 000--01010    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   212 | 11-0011010    | ...111.........1......1....1.1.. . . . . ...  . 1 1 .  . 1. .. .. .. . .  . . . .......... ... .      |
--   213 | 1--0011010    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   214 | --11011010    | .........11...11..............1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   215 | 01-1011010    | .1.............11....1........1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   216 | -0-0111010    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   217 | 1--0111010    | ................................ . . . . ...  . . 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   218 | 01-1111010    | .1111....1....1.....1111111..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   219 | 1-0-111010    | .1.1......1...1.1...........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   220 | 0-1-111010    | .1.1.1.........11..1..111.11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   221 | -010-11010    | ................................ . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   222 | 1001-11010    | 1..11....1....................1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   223 | 1101-11010    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   224 | 011--11010    | .1.1.1........1.1111111..111..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   225 | 00010-1010    | ...............................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   226 | -0101-1010    | 1..11....1...................... . . . . ...  . 1 . 1  . .. .. .1 .1 1 .  . . . .......... ... .      |
--   227 | 10-01-1010    | .1.1.1...1....1.11........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   228 | 000100-010    | ..111..........................1 . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   229 | 01-100-010    | .1111.....1...1......11111...11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   230 | 101--0-010    | ..111..........................1 . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   231 | 000001-010    | ................................ . . . . ...  . 1 . .  . .. 11 .. .. . .  . . . .......... ... .      |
--   232 | 010001-010    | ..1111...1....1..1.1.1.1.1.1.1.1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   233 | 1-1-01-010    | 1..111....................11..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   234 | --1011-010    | ................................ . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   235 | 01-011-010    | ..1111....1....1.1.1.1.1.1.1.1.1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   236 | 0--1-1-010    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... 1.. .      |
--   237 | 11-0000110    | 1...1.....1..................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   238 | 0001000110    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   239 | 1101000110    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   240 | --11000110    | ..111....11...11...........1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   241 | 10-1000110    | .1...1....1.............1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   242 | 11-1000110    | 1..11....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   243 | 011-000110    | .1...1.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   244 | 0000100110    | ...1.1...1...........111..11.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   245 | 0-01100110    | ..111..........................1 . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   246 | 0000-00110    | ................................ . . . . ...  . . . .  . .. 1. .. .. . .  . . . .......... ... .      |
--   247 | -010-00110    | ................................ . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   248 | 10-1-00110    | ................................ . . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   249 | 01-1-00110    | .11111...1................111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   250 | 11-0010110    | .1.1......1...1.11..........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   251 | 0001010110    | ..111.....1.....11111111111111.1 . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   252 | 0-11010110    | .11111.............1......11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   253 | -000110110    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   254 | 110-110110    | .11111....1..........1.11.111.1. . . . . ...  . . . .  . .. .. 1. .. . .  . . . .......... ... .      |
--   255 | 1001-10110    | 1..11....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   256 | 1101-10110    | .11111....1..........1.11111111. . . . . ...  . . . .  . .. .. 1. .. . .  . . . .......... ... .      |
--   257 | 011--10110    | .1111....1....1.....1111111..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   258 | 1-1-0-0110    | .........1.........11...1....... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   259 | 01001-0110    | .1.1.1........11111....1..11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   260 | 10011-0110    | .1...1...1.............11.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   261 | 0-111-0110    | .1.1.1....1...1.1....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   262 | 01-11-0110    | .1111...........11...11...1..... . . . . ...  1 . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   263 | 10-1--0110    | ................................ . . . . ...  . 1 . 1  . .. .. .. .. . .  . . . .......... ... .      |
--   264 | 0100001110    | .1.1.1........11111....1..11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   265 | -010001110    | ................................ . . . . ...  1 . . .  . .. .1 .1 .1 1 1  . . . .......... ... .      |
--   266 | 11-0001110    | ...111....................111... . . . . ...  1 . . .  . 11 .. .1 .. . .  . . . .......... ... .      |
--   267 | 0-11001110    | .1.1.1....1...1.1....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   268 | 01-1001110    | .11111.............1......111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   269 | 0000101110    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   270 | 10-0101110    | .1.1......1...1..1...1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   271 | 0-11101110    | ...1.1....1...11...1..1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   272 | 11--101110    | ...11....1....1.11............1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   273 | 1101-01110    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   274 | 011--01110    | .1...1...11...1...........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   275 | 11-0011110    | .1111....1....1..1...1.1111..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   276 | --11011110    | .....1....1....1........11.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   277 | -01-011110    | ................................ . . . . ...  1 1 . .  . .. .. .1 .. . .  . . . .......... ... 1      |
--   278 | -1-1111110    | .1.1.1........1.1111111..111..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   279 | -0--111110    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   280 | 11--111110    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   281 | 0000-11110    | ..........1.....11111111111111.. . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   282 | -010-11110    | .1...1...1.............11.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   283 | 0001-11110    | .1.......1....1.11............1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   284 | 10-1-11110    | .1.1.1........1..1........1111.. . . . . ...  1 . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   285 | 11-1-11110    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   286 | 00011-1110    | ................................ . . . . ...  . 1 . .  . .. 11 .. .. . .  . . . .......... ... .      |
--   287 | 00-11-1110    | .11.1....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   288 | 1--11-1110    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   289 | 01-110-110    | .1111.....1....1..11111...1..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   290 | 111-10-110    | 1..111........11........111111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   291 | --10-0-110    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   292 | 000001-110    | 1...1..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   293 | 0-1011-110    | .1...1...1.............11.1.111. . . . . ...  . 1 . 1  . .. .. .1 .. . .  . . . .......... ... 1      |
--   294 | 01-011-110    | .11111...1.....1...11.....111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   295 | -00111-110    | .1.1..........1......11...11111. . . . . ...  . . 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   296 | 110--1-110    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   297 | 11011--110    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   298 | -1111--110    | ................................ . . . . ...  . 1 . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   299 | 101----110    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   300 | -010000-10    | ................................ . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   301 | 01-1100-10    | .1.1.1.........111....1...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   302 | 0-00110-10    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   303 | 10-0110-10    | .1.1.1...1....1..1........1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   304 | 100-110-10    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   305 | --101-0-10    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   306 | 0000001-10    | .1...1.............11...1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   307 | 000-001-10    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   308 | 11-0101-10    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   309 | 111-101-10    | 1..111...1....11........111111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   310 | 0000011-10    | .....1...............111..11.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   311 | 00--011-10    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   312 | -001111-10    | ...............................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   313 | 101--11-10    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   314 | 00010-1-10    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   315 | 1-0-1-1-10    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . 11..111... 1.. .      |
--   316 | -0-100--10    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . 1..1..11.1 ... .      |
--   317 | 01-1-0--10    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   318 | 1-0111--10    | ...111...1.............11.1.111. . . . . ...  . . . 1  . .. .. .1 .. . .  . . 1 .......... ... .      |
--   319 | 00000---10    | .........1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   320 | 1--00000-0    | ................................ . . . . ...  . . . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   321 | -0101000-0    | .1.......1....1.11............1. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   322 | 10-10100-0    | ..111........................1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   323 | 01-10100-0    | .11111.............11.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   324 | -01-0100-0    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   325 | 11-00-00-0    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   326 | -0-00010-0    | .................1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   327 | 11-00010-0    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   328 | 000-0010-0    | .1.1......1...1.11..........111. . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   329 | 0000-010-0    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   330 | 01-0-010-0    | ................................ . . . . ...  . 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   331 | 1--00110-0    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   332 | 0-010110-0    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   333 | -0-1-110-0    | ................................ . . . . ...  1 . 1 1  . .. .. .. .. . .  . . . .......... ... .      |
--   334 | 10-000-0-0    | ................................ . . . . ...  . . . .  . .1 .. .1 .. . .  . . . .......... ... .      |
--   335 | 1-1-0001-0    | 1..111....1..............1111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   336 | 11--0001-0    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   337 | 10-01001-0    | ..111........................1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   338 | 01-11001-0    | ..111....1.....................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   339 | 10-1-001-0    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   340 | -0100101-0    | .................1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   341 | 11-00101-0    | ................................ . . . . ...  . . 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   342 | 11-0-011-0    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   343 | 10-1-111-0    | ..............................1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   344 | 101--111-0    | ...111.............1.1..11111... . . . . ...  . . 1 .  . .1 .. .. .. . .  . . . .......... ... .      |
--   345 | 0-101-11-0    | .1.......1....1.11............1. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   346 | -1111-11-0    | 1..111.........1..........1...1. . . . . ...  . 1 1 1  . .1 .. .. .. . 1  . . . .......... ... .      |
--   347 | 000111-1-0    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   348 | 1-0111-1-0    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   349 | 10-01--1-0    | ................................ . . . . ...  1 . . .  . .. .. .. .. . .  . . 1 1...1..1.1 ... .      |
--   350 | 011-1--1-0    | .11111.........1....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   351 | 10-0000--0    | 1............................... . . . . ...  . . . .  . .1 .1 .1 .1 1 1  . . . .......... ... .      |
--   352 | 11-0100--0    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   353 | -110110--0    | 1....1...1................1..... . . . . ...  1 . . .  . .. .. 11 .. . .  . . . .......... ... .      |
--   354 | 0000001--0    | ................................ . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... 1      |
--   355 | 10--001--0    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   356 | 1-1-011--0    | 1...11.........1..........1...1. . . . . ...  . . 1 .  . .1 .. .. .. . 1  . . . .......... ... .      |
--   357 | -001111--0    | 1..11....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   358 | 10-00-1--0    | ....1........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   359 | 0001000001    | 1...1....1...................... . . . . ...  . . . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   360 | 0-11000001    | ...............11....1.......... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   361 | 110-000001    | .1.1.1....1...1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   362 | 011-000001    | .1111....1....1.....1111111..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   363 | 0-11100001    | .11111...11...1.........11.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   364 | 1-1-100001    | 1....1....1...............11..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   365 | 0000-00001    | 1...1.....1..................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   366 | 11-0-00001    | .1111....1....1.11............1. . . 1 . ...  . . . .  . .. .. .. .. . .  . 1 . .......... 1.. .      |
--   367 | 000-010001    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   368 | 010-010001    | .1111.........111....1........1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   369 | -000110001    | ................................ . . . . ...  . 1 1 .  . .. 11 .. .. . .  . . . 1...1.1..1 ... .      |
--   370 | -1-0110001    | .11.1.....1...1................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   371 | 00-1110001    | .1.1.1....1...1.1....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   372 | -00-110001    | ................................ . 1 . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   373 | -11-110001    | 1..111....................11..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   374 | 1101-10001    | .11111...1.............11.1.111. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   375 | 10-1-10001    | ................................ . . . . ...  . . 1 .  . .1 .. .. .. . .  . . . .......... ... .      |
--   376 | 011--10001    | .11111....1....1...1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   377 | 1-1--10001    | .........1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   378 | 01000-0001    | ..111....1.......1.1.1.1.1.1.1.1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   379 | 11-00-0001    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   380 | --010-0001    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . ......11.. ... .      |
--   381 | 1-1-0-0001    | 1..111....1...............1111.. . . . . ...  1 . 1 1  . .. 1. .. .. . .  . . . .......... ... .      |
--   382 | 01001-0001    | .11111...1.....1...11.....111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   383 | 10011-0001    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   384 | 11011-0001    | ................................ 1 . . . ...  . . . .  . 1. .1 .1 .1 1 1  . . . .......... ... .      |
--   385 | 101---0001    | ...................1.1..11...... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   386 | 0-00001001    | .11111...1.....1...11.....111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   387 | --10001001    | .1111....1....1....11111..1..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   388 | 11-1001001    | 1..11....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   389 | ---1001001    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   390 | -01-001001    | .1.1.1....1...1.1....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   391 | -000101001    | 1...1....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   392 | 0100101001    | .1.1.1........1111....1...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   393 | 11-0101001    | ..111...................1....11. . . . . ...  . . 1 .  . .. .1 .. .. . .  . . . .......... ... 1      |
--   394 | 0001101001    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   395 | 0-11101001    | ..111....11...11...........1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   396 | 01-1101001    | .1.1.1........1.1111111..111..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   397 | 11-1101001    | ................................ . . . . ...  1 1 . 1  . .. .. .1 .. . .  . . . .......... 1.. 1      |
--   398 | 11-0011001    | ..111.....1.....11111111111111.1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   399 | 0001011001    | 1...1....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   400 | 01-1111001    | .11111...11...1...........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   401 | 1-0-111001    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   402 | 0000-11001    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   403 | --10-11001    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   404 | 1101-11001    | .1111.....1....1.1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   405 | 0-11-11001    | .11111.............1......11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   406 | 101--11001    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   407 | 10-01-1001    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   408 | 11011-1001    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   409 | 1-011-1001    | .11111...1.............11.1.111. . . . . ...  . . . 1  . .. .. .1 .. . .  . . . .......... ... .      |
--   410 | 00--1-1001    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . ....1..11. ... .      |
--   411 | -01000-001    | .1.1..........1......11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   412 | 11-000-001    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   413 | 01-100-001    | .....1.........1................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   414 | -00-10-001    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . ...1...11. ... .      |
--   415 | 101--0-001    | .11111...1..............1.1.111. . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   416 | 010001-001    | ..111....1.......1.1.1.1.1.1.1.1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   417 | 0-1101-001    | .11111.............1......11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   418 | 0-1011-001    | .1111.....1...1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   419 | 01-011-001    | ..111.....1......1.1.1.1.1.1.1.1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   420 | 1101000101    | ................................ . . . . ...  1 . . .  . .. .1 .1 .1 1 1  . . . .......... ... .      |
--   421 | 10-1000101    | .1.1......1...1..1...1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   422 | 01-1000101    | .11111...1.....1...11.....111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   423 | 000-000101    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   424 | 011-000101    | .1.1.1........1.1111111..111..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   425 | 1-1-000101    | 1..111..................1.1111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   426 | 11-0100101    | .11111.............1.1..1111111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   427 | 1--0100101    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   428 | 0001100101    | .1...1..................1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   429 | 0-01100101    | ................................ . . . . ...  . . 1 .  . .. .1 .. .. . .  . . . .......... ... 1      |
--   430 | 0-11100101    | .1...1.........1........11.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   431 | 1-1-100101    | 1....1...1.....1....1.....111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   432 | 10--100101    | ................................ . . 1 . ...  . . . .  . .1 .. .. .. . .  . . 1 .......... ... .      |
--   433 | 11-0010101    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   434 | 0001010101    | .11111...1...........1111.11.1.. . . . . ...  . . . .  . .. 11 .. .. . .  . . . .......... ... .      |
--   435 | -101010101    | .11111.............11.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   436 | -01-010101    | .11111...11...11...1..1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   437 | 0-00110101    | ...1....................1.1.111. . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... 1      |
--   438 | 110-110101    | .11111.........1......1....1.1.. 1 . . . ...  . 1 1 .  . 1. .. .. .. . .  . . . .......... ... .      |
--   439 | 01--110101    | ..........1....1................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   440 | 1101-10101    | ................................ 1 . . . ...  . . . .  . 1. .1 .. .. . .  . . . .......... ... .      |
--   441 | 011--10101    | .11111...11...1...........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   442 | 01000-0101    | .11111.........1.........1.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   443 | -0100-0101    | .11111...1.............11.1.111. . . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... 1      |
--   444 | 1-1-0-0101    | ................................ . . . . ...  . . . .  . .. 1. 11 .. . .  . . . .......... ... .      |
--   445 | 0-001-0101    | .....1........1................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   446 | 0-111-0101    | ..111.....1.....11.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   447 | -1-11-0101    | ................................ . . . . ...  . 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   448 | 101---0101    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   449 | 0100001101    | .....1........1................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   450 | 11-0001101    | ................................ 1 . . . ...  . . . .  . 1. .1 .1 .1 1 1  . . . .......... ... .      |
--   451 | 0001001101    | .11111...1..............1.1.111. . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   452 | 01-1001101    | .11111.............11.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   453 | 0-11101101    | .1.1.1...1....1......111..111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   454 | 01-1101101    | .1111.....1....1....1111111..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   455 | -010-01101    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   456 | 11-0-01101    | ..111.........1.....1.11.1.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   457 | 10-1-01101    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . 1 1.111.1.1. ... .      |
--   458 | 011--01101    | .11111.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   459 | --11011101    | ...............1..........1...1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   460 | 11--011101    | ................................ . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   461 | -1-1111101    | .1111................11...1...1. . . . . ...  1 . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   462 | 0000-11101    | ................................ . . . . ...  . 1 . .  . .. 11 .. .. . .  . . . .......... ... .      |
--   463 | 11-0-11101    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   464 | 0001-11101    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   465 | 1001-11101    | ..111........................1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   466 | -0-1-11101    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   467 | 11-1-11101    | 1..11....1...................... . . . . ...  . . . 1  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   468 | 0-1100-101    | ..111.....1.....1111............ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   469 | 000010-101    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   470 | --0010-101    | ................................ . . . . ...  . 1 1 .  . .. .. .. .. . .  . . . ....1.1.1. ... .      |
--   471 | 000110-101    | ..111....1.....1................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   472 | 101--0-101    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   473 | -00001-101    | 1...1.....1..................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   474 | 010001-101    | .11111.........1.........1.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   475 | -01001-101    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   476 | 01-011-101    | .1111.........1111111....1....1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   477 | 11011--101    | .1........1....1.1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   478 | 011-1--101    | .1.1.1....1.....11....1...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   479 | 11-0000-01    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   480 | -010100-01    | .1111.....1...1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   481 | 10-1100-01    | .1.1.1........1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   482 | -010010-01    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   483 | 10-1010-01    | ................................ . . 1 . ...  1 . . .  . .1 .. .. .. . .  . . 1 .......... ... .      |
--   484 | 10-0110-01    | ...1.1........1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   485 | 0001110-01    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . 1 . .......... ... .      |
--   486 | 01--110-01    | .11111.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   487 | 1101-10-01    | ................................ . . . . ...  . . . 1  . .. .. .1 .. . .  . . . .......... ... .      |
--   488 | -01--10-01    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . ........1. ... .      |
--   489 | 0000001-01    | ..111....11....................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   490 | 10-1001-01    | .1.1.1...1....1..1........1.111. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   491 | 11-0101-01    | .1...1...1................1.1... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   492 | -1-0-01-01    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   493 | 01---01-01    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   494 | -001111-01    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   495 | 100-111-01    | ...1.1..................1.1.111. . . 1 . ...  . 1 . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   496 | 011--11-01    | .1111................11...1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   497 | -0101-1-01    | .1111....1....1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   498 | -00011--01    | .11.1....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   499 | 00000---01    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   500 | 0-------01    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   501 | -010000011    | .1...1...1.............11.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   502 | 1101000011    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   503 | 011-000011    | .11111....1....1...1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   504 | 1-1-000011    | .........11.........1....1..1... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   505 | -010100011    | .1111.....1....1.1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   506 | 1--0100011    | .1.1.....1.....1.....11...11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   507 | 0-11100011    | .11111.............1.1....11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   508 | 0000-00011    | .1.1......1...1..1...1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   509 | 10-1-00011    | .1...1....1.............1.1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   510 | 10---00011    | ................................ . . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   511 | -000010011    | .....1................1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   512 | -010010011    | ................................ . . . . ...  . . . .  . 1. .. .. .1 1 .  . . . .......... ... .      |
--   513 | -0-0010011    | ..111........................... 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   514 | 1--0010011    | .11111...1....1.....1.11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   515 | 10--010011    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   516 | -101110011    | .........1..........11111.1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   517 | 00-1110011    | .11111...11...11...1..1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   518 | 0-00-10011    | ................................ . . . . ...  . . 1 .  . 1. .1 .. .. . .  . . . .......... ... .      |
--   519 | 0001-10011    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   520 | 1101-10011    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   521 | 011--10011    | .1.1.1........1.1111111..111..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   522 | 01000-0011    | .1.1.1........1111111....111111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   523 | -0100-0011    | ................................ . . . . ...  . . . .  . .. .1 .1 .. . .  . . . .......... ... 1      |
--   524 | 0-110-0011    | .1.1.1....1...1.1....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   525 | ---10-0011    | ................................ . . . . ...  1 . . .  . .. .. .. .. . .  . . . .1.......1 ... .      |
--   526 | -11-0-0011    | ................................ . . . . ...  . 1 1 1  . .. .. .. .. . .  . . . .......... ... .      |
--   527 | 10-01-0011    | 1...1.....1..................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   528 | 00011-0011    | ................................ 1 . . . ...  . . . .  . 1. .1 .1 .1 1 .  . . . .......... ... .      |
--   529 | 101---0011    | ................................ . . . . ...  1 . . .  . 11 .. .1 .. . .  . . . .......... ... .      |
--   530 | 1--0001011    | .1...1.............1.1..111111.. . . . . ...  . . 1 .  . .1 .. .. .. . .  . . . .......... ... .      |
--   531 | 1101001011    | .1...1....1..........1.1111111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   532 | 00-1001011    | .11111...11...11...1..1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   533 | 11-1001011    | ................................ . . . . ...  1 . . .  . .. .. 1. .. . .  . . . .......... ... .      |
--   534 | 0000101011    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   535 | 11-0101011    | .1.......1....1..1...1.1111..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   536 | 01-1101011    | .1............11................ . . . . ...  1 . . .  . 11 .. .. .. . .  . . . .......... ... .      |
--   537 | 0-1-101011    | ..111.....1.....11111111........ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   538 | 0001-01011    | .1........1....1.1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   539 | 011--01011    | .1111...........1....11...1...1. . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   540 | 1--0011011    | ................................ . . . . ...  . . . .  . .. .. .1 .1 1 1  . . . .......... ... .      |
--   541 | --11011011    | .11111........1....11....1.1.... 1 . . . ...  . . . .  . 1. .. .. .. . 1  . . . .......... ... .      |
--   542 | 0---011011    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   543 | -1-1111011    | .1.......1....1...1.111.1.1..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   544 | -010-11011    | .11111...1.............11.1.111. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   545 | 11-0-11011    | ................................ . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   546 | 11-1-11011    | .1........1...1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   547 | 00010-1011    | .1111....1....1..1...1.1111..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   548 | --101-1011    | ................................ 1 . . . ...  . . . .  . 1. .1 .1 .1 1 .  . . . .......... ... .      |
--   549 | 11----1011    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   550 | 000100-011    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   551 | 01-100-011    | .11111....1...1....1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   552 | 10-110-011    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   553 | -00001-011    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   554 | 010001-011    | .1.1.1........1111111....111111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   555 | 1-1-01-011    | 1...11....1.............11111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   556 | 000011-011    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   557 | --1011-011    | .11111...1.............11.1.111. . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   558 | 01-011-011    | .1111.....1...1......11111...11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   559 | 000111-011    | ................................ 1 . . . ...  . . . .  . 1. .1 .1 .1 1 1  . . . .......... ... .      |
--   560 | -010-1-011    | ................................ . . . . ...  . . . .  . .. .. .1 .. . 1  . . . .......... ... 1      |
--   561 | 0-011--011    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   562 | 011-1--011    | .1.1.1....1.....111....1..11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   563 | 111-1--011    | 1..111.........1....1...1.1111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   564 | -1-1---011    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   565 | --00000111    | ..............1................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   566 | -010000111    | .11111................1....1.1.. . . . . ...  . . . .  . 1. .. .1 .. . .  . . . .......... ... .      |
--   567 | -0-0000111    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   568 | 0001000111    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   569 | 0-11000111    | .11111.............1.1....11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   570 | 011-000111    | .11111...11...1...........11.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   571 | -010100111    | 1..11....1...................... . . 1 . ...  . . . .  . .. .. .1 .1 1 .  . . . .......... ... .      |
--   572 | 11-0100111    | ................................ . . . . ...  . . . .  . 1. .1 .1 .1 1 1  . . . .......... ... .      |
--   573 | 1--0100111    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   574 | 0-01100111    | .1111....1....1..1...1.1111..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   575 | 0-11100111    | .1.1.1...1....1......11.1111.11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   576 | -000-00111    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   577 | 11-0-00111    | ..111...............1.11.1.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   578 | 0-00010111    | .1.1......1...1..1...1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   579 | 1--0010111    | .11111.............1.1..111111.. . . . . ...  . . 1 .  . .1 .. .. .. . .  . . . .......... ... .      |
--   580 | 0-01010111    | .11111.........1......1....1.1.. 1 . . . ...  . . . .  . 1. .. .. .. . .  . . . .......... ... .      |
--   581 | 0-11010111    | .1.1.1.........11..1..111.11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   582 | 110-110111    | .1.1.1....1...1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   583 | 010--10111    | .1.1.1..........1111111...11..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   584 | 01-10-0111    | .11111..............1.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   585 | -000001111    | .1.1......1...1..1...1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   586 | -010001111    | 1..11....1...................... . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   587 | 1--0001111    | ..111...................1....11. . . . . ...  1 . 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   588 | --11001111    | .1.1.1...1....1......111.1111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   589 | 10--001111    | .11.1....1...................... 1 . . . ...  . 1 . .  . .. 11 .. .. . .  . . . .......... ... .      |
--   590 | 0-00101111    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   591 | 0001101111    | ..111.....1.....1111111111111..1 . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   592 | -1-1101111    | ................................ . . . . ...  1 . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   593 | 11--101111    | .1111.....1....1.1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   594 | 0--0-01111    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   595 | 11-1-01111    | .1.1......1...1.1...........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   596 | -0-0011111    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   597 | 1--0011111    | 1...1.....1..................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   598 | 0-01011111    | .1111.....1....1.1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   599 | 00-0111111    | .11111.........1......1....1.1.. 1 . . . ...  . 1 1 .  . 1. .. .. .. . .  . . . .......... ... .      |
--   600 | 11--111111    | .11111...1.............11.1.111. 1 . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   601 | --10-11111    | .1...1................1....1.1.. 1 . . . ...  . . . .  . 1. .1 .1 .. . .  . . . .......... ... .      |
--   602 | 10-0-11111    | .1.1.1...1....1.11........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   603 | --11-11111    | ..........1...1...........1...1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   604 | 10-1-11111    | 1..11....1...................... . . 1 . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   605 | 01-1-11111    | .11111.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   606 | 11-1-11111    | .1111....1....1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   607 | 01-10-1111    | .1111.........1111....1.......1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   608 | --101-1111    | .1111.....1....1.1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   609 | 1-011-1111    | .11111...1.............11.1.111. . . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   610 | 0-111-1111    | .11111.............1......11.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   611 | -11---1111    | .1111....1....1.....1111111..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   612 | 1-1---1111    | .1.1.....1....1.1....1....1.111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   613 | 11-000-111    | .1...1...1................1.1... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   614 | 01-110-111    | .1111...........1....11...1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   615 | 111-10-111    | 1....1....1........11...1.111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   616 | 0100-0-111    | .....1.............1............ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   617 | 010-01-111    | .....1........1................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   618 | 0-1011-111    | ................................ . . . . ...  . . . .  . 1. .1 .1 .. . .  . . . .......... ... .      |
--   619 | --1011-111    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   620 | 01-011-111    | .11111.........1.........1.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   621 | 0-1111-111    | .1.1.....1....1......1.11.1.1... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   622 | 0-1-11-111    | .....1................1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   623 | 1-01-1-111    | ................................ . . . . ...  1 1 . 1  . .. .. .. .. . .  . . . 11.1.111.1 ... .      |
--   624 | 101--1-111    | .11111....1.............1.1.111. . . . . ...  . . 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   625 | 011--1-111    | .1111....1....1.....11111.1..1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   626 | 011-1--111    | .1.1.1....1.....1....1....11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   627 | -10-000-11    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . 11.....1.. ... .      |
--   628 | ----100-11    | ................................ . . . . ...  . . 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   629 | 010-010-11    | ..111.....1..............1111111 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   630 | 0-00110-11    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   631 | 0001110-11    | ................................ . . . . ...  . . . .  . .. .1 .1 .1 1 1  . . . .......... ... .      |
--   632 | -001110-11    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   633 | -1-1110-11    | ..............1..........1...... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   634 | 01001-0-11    | .11111..............1.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   635 | 11011-0-11    | .1........1...1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   636 | 01--1-0-11    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   637 | -1-0--0-11    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   638 | 0100001-11    | .11111..............1.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   639 | 0001001-11    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   640 | 01-0101-11    | ..111....1................111111 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   641 | 10-0-01-11    | ....1.....1....................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   642 | 0-1-111-11    | .1.1.1....1...1.11111....111111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   643 | -11--11-11    | .11111.............1..11.1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   644 | 1-1--11-11    | .1.1......1...1.11..........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   645 | 0-010-1-11    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   646 | -1110-1-11    | .........1..............1....... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   647 | 11011-1-11    | .1.......1....1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   648 | -1-1--1-11    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   649 | 11-111--11    | ................................ . . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   650 | -1--11--11    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   651 | 1-10----11    | ................................ . . . . ...  . 1 1 .  1 .1 .. .. .1 1 1  . . . .......... ... .      |
--   652 | 11-00000-1    | 1...1....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   653 | 10--0000-1    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   654 | 01-11000-1    | .1...1....1...........1..1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   655 | ---11000-1    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   656 | -1-00100-1    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . 11...1.... ... .      |
--   657 | 10-10100-1    | 1..1............................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   658 | 10--0100-1    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   659 | 00011-00-1    | ..111....1.....1................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   660 | 101---00-1    | .11111....................111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   661 | -0000010-1    | ................................ . . . . ...  . . . .  . 1. .. .1 .. . .  . . . .......... ... .      |
--   662 | -0100010-1    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   663 | 00010010-1    | .11111...1...........1111.11.1.. 1 . . . ...  . . . .  . .. 11 .. .. . .  . . . .......... ... .      |
--   664 | 111-1010-1    | 1..111.........1.........11111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   665 | 11-00110-1    | ................................ . . . . ...  1 . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   666 | 1001-110-1    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   667 | 101--110-1    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   668 | 10-000-0-1    | ..111........................... 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   669 | 0-1-11-0-1    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   670 | -0-10--0-1    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   671 | 1001---0-1    | ................................ . . . . ...  1 . . .  . .. .. .. .. . .  . . 1 1....11..1 ... .      |
--   672 | 11010001-1    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   673 | --1-0001-1    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   674 | 01-11001-1    | .1...1.............1......111... 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   675 | 0--0-001-1    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   676 | -0100101-1    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   677 | 10-10101-1    | .1.1.1...1....1..1........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   678 | 100-1101-1    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   679 | 1-0-1101-1    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   680 | 1101-101-1    | .1111.....1...1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   681 | 0--10-01-1    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   682 | 11010011-1    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   683 | 10-01011-1    | ....1.....1...................1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   684 | 01-01011-1    | .11111.............11.1....1.1.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   685 | 10-00111-1    | .11...........................1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   686 | -1--0111-1    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... 1.. .      |
--   687 | ---01111-1    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   688 | 1--11111-1    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   689 | 0-1-1111-1    | ..111....11...11..............1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   690 | -11--111-1    | .........1....1.....1..111...... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   691 | 10-00-11-1    | 1...1........................... . . . . ...  . 1 . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   692 | -1110-11-1    | 1..111.........1..........1...1. . . . . ...  . 1 1 1  . .1 .. .. .. . 1  . . . .......... ... .      |
--   693 | 11011-11-1    | .....1................1....1.1.. . . . . ...  . . . .  . 1. .1 .1 .. . .  . . . .......... ... .      |
--   694 | 11-11-11-1    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   695 | ----00-1-1    | ................................ . . . . ..1  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   696 | 1-1--0-1-1    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   697 | 1-1-01-1-1    | 1...11...................11111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   698 | 0-1011-1-1    | .1111....1....1..1.............. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   699 | 1-0111-1-1    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   700 | 11-111-1-1    | .........1..............1....... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   701 | 0-11---1-1    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   702 | 10-0000--1    | ...11........................... 1 . . . ...  . . . .  . 1. .1 .1 .1 1 1  . . . .......... ... .      |
--   703 | 10-0100--1    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   704 | -1-1100--1    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   705 | 10-00-0--1    | ..1............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   706 | 00-10-0--1    | ................................ . . . . ...  . 1 1 .  . .. .. .. .. . .  . . . ...1....1. ... .      |
--   707 | -1111-0--1    | ................................ . . . . ...  1 1 . 1  . .. .. .. .. . .  . . . .......... ... .      |
--   708 | 01-1011--1    | .11111....1...........1..1111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   709 | 1-1-011--1    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   710 | 11-1111--1    | ................................ . . . . ...  . 1 1 1  . .1 .. .. .. . 1  . . . .......... ... .      |
--   711 | -11-111--1    | 1...11.........1..........1...1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   712 | 1-001-1--1    | ................................ . . . . ...  1 . . .  . .. .. .. .. . .  . . 1 11........ ... .      |
--   713 | 011-1-1--1    | .11111....1............1..1..... . . . . ...  . . . .  . .. .1 .1 .. . .  1 . . .......... ... .      |
--   714 | 1-10--1--1    | ................................ 1 . . . ...  . . 1 .  1 .1 .1 .. .1 1 1  . . . .......... ... .      |
--   715 | 10-010---1    | 1............................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   716 | 10-001---1    | 1............................... . . . . ...  . 1 . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   717 | 0-1-1----1    | ................................ . . . . ...  . . . 1  . .. .. .. .. . .  . . . ..1.1....1 1.. .      |
--   718 | 1-10-----1    | 1..111....1...1.....1.....1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   719 | 0-1100000-    | .1.1.1....................11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   720 | 01-100000-    | ..111.....1.......11..11..11..11 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   721 | -1-010000-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . 11...111.1 ... .      |
--   722 | 000110000-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . ...1.1111. ... .      |
--   723 | 01-110000-    | ................................ . . . . ...  1 . 1 .  . .1 .. .. .. . .  . . . .......... ... .      |
--   724 | -010-0000-    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   725 | 1--11-000-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   726 | 011-1-000-    | .1.1.1.........1.............11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   727 | -0-000100-    | ................................ . . . . ...  . . . .  . .. .1 .. .1 1 .  . . . .......... ... .      |
--   728 | 01-100100-    | ..111.....1.........1111....1111 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   729 | 1-1-00100-    | 1..111....1........1....11111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   730 | 11--00100-    | ................................ . . . . ...  1 1 1 1  . .. .. .. .. . .  . . . 11.1...11. ... .      |
--   731 | 0-1101100-    | ..........1...1..........1..1... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   732 | 01-101100-    | ................................ . . . . ...  . . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   733 | 100-11100-    | .11.1....1...................... 1 . . . ...  . 1 . .  . .. 1. .. .. . .  . . . .......... ... .      |
--   734 | 1--0-1100-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   735 | 0----1100-    | ................................ . . . . ...  1 . 1 .  . .. .. .. .. . .  . . . .....1.... ... .      |
--   736 | -0100-100-    | .1.1..........1.1...........111. . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   737 | -01000-00-    | ................................ . . . . ...  . . 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   738 | 11-000-00-    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   739 | 000001-00-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   740 | 0-1011-00-    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . ..1.1.111. ... .      |
--   741 | 0--111-00-    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   742 | 110-11-00-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . 11..1.111. ... .      |
--   743 | --1-11-00-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   744 | ---0---00-    | ................................ . . . . 1.1  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   745 | 0-1100010-    | .1...1...1....1.........11.1.... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   746 | 0-0-00010-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   747 | 00-010010-    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . ..1.1...1. ... .      |
--   748 | 0000-0010-    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   749 | 11-001010-    | ................................ . . . . ...  . . 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   750 | -1-1-1010-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   751 | 01001-010-    | ..111....1..........1111....1111 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   752 | 101---010-    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   753 | 010000110-    | ..111....1..........1111....1111 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   754 | 1--000110-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   755 | 110100110-    | .1.1.1....1...1...........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   756 | 0-0-01110-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . ...1.11.1. ... .      |
--   757 | -100-1110-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   758 | 00011-110-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   759 | 10011-110-    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   760 | 10-100-10-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . 1..1..1..1 ... .      |
--   761 | ----01-10-    | ................................ . . . . 1.1  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   762 | 000111-10-    | .1.1.1........1.1...........111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   763 | 11-111-10-    | 1...11....1........11...1.111.1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   764 | 0-10-1-10-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .....1.... ... .      |
--   765 | 0-1-010-0-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......1.. ... .      |
--   766 | -110110-0-    | ................................ . . . . ...  1 . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   767 | 01-1-10-0-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   768 | 11-00-0-0-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   769 | 0-0-1-0-0-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   770 | -010001-0-    | .1.1..........1.1...........111. . . . . ...  . . 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   771 | 1001-11-0-    | ................................ . . . . ...  1 1 . 1  . .. .. .. .. . .  . . . 1..1.1.1.1 ... .      |
--   772 | 0--0-0--0-    | ................................ . . . . ...  1 . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   773 | --0111--0-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   774 | -01000001-    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   775 | 110100001-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   776 | -01010001-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . 1 . .......... 1.1 .      |
--   777 | 11-010001-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . 1 . 11..1....1 ... .      |
--   778 | 10--10001-    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   779 | 0-00-0001-    | ................................ . . . . ...  . 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   780 | 10-0-0001-    | ................................ . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   781 | -0-1-0001-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   782 | -0-001001-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   783 | -0--01001-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   784 | 000-11001-    | ................................ 1 . . . ...  . . . .  . 1. .1 .1 .1 1 1  . . . .......... ... .      |
--   785 | -1--11001-    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   786 | 0001-1001-    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   787 | -00100101-    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   788 | 0001-0101-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . 1 . .......... 1.. .      |
--   789 | 00-011101-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   790 | 100-11101-    | ..111....1...................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   791 | 01---1101-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   792 | 1-1-0-101-    | 1..111...................11111.. . . . . ...  1 . . 1  . .. 1. 11 .. . .  . . . .......... ... .      |
--   793 | -1--0-101-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   794 | --1-1-101-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   795 | -00001-01-    | .11.1........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   796 | 0-0001-01-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   797 | ---111-01-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   798 | 1-01-1-01-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . 1..1.1.... ... .      |
--   799 | 10-00--01-    | ..1............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   800 | 000100011-    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   801 | 0000-0011-    | .11.1........................... . . . . ...  . 1 . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   802 | -000-0011-    | ................................ . 1 . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   803 | 10-1-0011-    | ..111..........................1 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   804 | ---1-0011-    | ................................ . . . . ...  1 1 . 1  . .. .. .. .. . .  . . . .......... ... .      |
--   805 | 010-01011-    | .11111..............1.....111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   806 | 0-00-1011-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   807 | 01000-011-    | ..111....1........11..11..11..11 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   808 | -1-01-011-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   809 | -1--1-011-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   810 | 1---00111-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   811 | 00-010111-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . 1 . .......... 1.1 .      |
--   812 | 01-010111-    | .11111.............1......111... 1 . . . ...  . 1 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   813 | ---110111-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   814 | 11--10111-    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   815 | 1101-0111-    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   816 | 000101111-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . 1 . .......... 1.. .      |
--   817 | 01-101111-    | .1111................111111..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   818 | --1-11111-    | .....1........1....11....1.1.... 1 . . . ...  . . . .  . 1. .. .. .. . 1  . . . .......... ... .      |
--   819 | -11--1111-    | .11111....1........1..11.1111... 1 . . . ...  . . 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   820 | --1--1111-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   821 | -111--111-    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   822 | 101--0-11-    | ................................ . . . . ...  . . 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   823 | 010001-11-    | ..111....1........11..11..11..11 . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   824 | 01-101-11-    | ................................ 1 . . . ...  . 1 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   825 | 1-1-01-11-    | ................................ . . . . ...  . . . .  . .. 1. 11 .. . .  . . . .......... ... .      |
--   826 | 1-0-11-11-    | ................................ . . . . ...  1 1 . 1  . .. .. .. .. . .  . . . .......1.. ... .      |
--   827 | --1-11-11-    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   828 | ---0-1-11-    | ................................ . . . . ..1  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   829 | -111-1-11-    | 1...11.........1.........11111.. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   830 | 011----11-    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   831 | 1-1-000-1-    | 1..111.........1..........11..1. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   832 | 01--100-1-    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   833 | 10-0110-1-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   834 | 01-0--0-1-    | ................................ . . . . ...  1 . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   835 | 010-001-1-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   836 | 111-101-1-    | ................................ . . . . ...  . . . .  . .. .. .1 .. . .  . . . .......... ... .      |
--   837 | 1---101-1-    | ................................ . . . . ...  1 1 . 1  . .. .. .. .. . .  . . . 11.11.1..1 ... .      |
--   838 | -----01-1-    | ................................ . . . . .11  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   839 | -000011-1-    | ................................ . . . . ...  . . . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   840 | 11-1111-1-    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   841 | 01--111-1-    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   842 | 101--11-1-    | ................................ . . . . ...  . 1 1 .  . .. .. .. .. . .  . 1 . .......... ... .      |
--   843 | 10-00-1-1-    | ................................ 1 . . . ...  . 1 . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   844 | -1101-1-1-    | ................................ 1 . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   845 | 011-1-1-1-    | .11111...1.....1......111.1..11. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   846 | -00010--1-    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   847 | 10-001--1-    | .11.1........................... 1 . . . ...  . 1 . .  . .. .1 .. .. . .  . . . .......... ... .      |
--   848 | -1--11--1-    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   849 | 1-011---1-    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   850 | 0-11----1-    | ................................ . . . . ...  . 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   851 | 10-01000--    | .11.1........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   852 | -110-000--    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   853 | 00011100--    | .11111.........1......1....1.1.. 1 . . . ...  . . 1 .  . 1. .. .. .. . .  . . . .......... ... .      |
--   854 | 00000010--    | .11111....................111... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   855 | -0100010--    | .1.1.1........1...........11111. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   856 | 00-00010--    | ................................ . . . . ...  1 . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   857 | --101110--    | 1..111....1...............1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   858 | 1101-110--    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . .1....1... ... .      |
--   859 | 100110-0--    | ................................ . . . . ...  1 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   860 | 0-00-0-0--    | ................................ . . . . ...  1 . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   861 | -1--11-0--    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   862 | -0100101--    | .1.1.1........1...........11111. . . . . ...  1 . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   863 | 100-1101--    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . 1...11..1. ... .      |
--   864 | -0011-01--    | ................................ . . . . ...  1 . . .  . .. .. .. .. . .  . . . ...1...... 1.. .      |
--   865 | 11011-01--    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . 1 . 11.11..1.. ... .      |
--   866 | --11--01--    | ................................ . . . . ...  1 . . 1  . .. .. .. .. . .  . . . .......... ... .      |
--   867 | -1010011--    | ................................ . . . . ...  1 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   868 | 10-01011--    | ................................ . . . . ...  . 1 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   869 | --110111--    | .1111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   870 | -0011111--    | .1.1.1........1.11........11111. . . . . ...  1 . . .  . .1 .. .. .. . .  . . . .......... ... .      |
--   871 | 1--11111--    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   872 | -1101-11--    | 1...11....1...............1..... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   873 | -1-11-11--    | ................................ . 1 . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   874 | 0--11-11--    | ................................ . . . 1 ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   875 | ---110-1--    | ................................ . . . . 11.  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   876 | 0-0001-1--    | ................................ . . . . ...  1 . 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   877 | 0000100---    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   878 | 0100-10---    | .11111.............1......111... 1 . . . ...  . 1 1 .  . .. .1 .. .. . .  . . . .......... ... .      |
--   879 | ----0-0---    | ................................ . . . . 1..  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   880 | ----111---    | ................................ . . . . 11.  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   881 | 11011-1---    | ..111........................... . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   882 | ----00----    | ................................ . . . . .1.  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   883 | ---0-0----    | ................................ . . . . 1..  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   884 | 0-11-0----    | ................................ . . . . ...  1 . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   885 | 011--0----    | ................................ . . . . ...  1 . 1 .  . .. .. .. .. . .  . . . .......... ... .      |
--   886 | ---111----    | ................................ . . . . .1.  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   887 | 0--00-----    | ................................ . . . . ...  . . . 1  . .. .. .. .. . .  . . . ..1...1.11 ... .      |
--   888 | 0-111-----    | ................................ . . . . ...  . 1 . .  . .. .. .. .. . .  . . . .......... ... .      |
--   889 | 111-------    | .11............................. . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   890 | --1-------    | ................................ . . . . 1.1  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   891 | -1--------    | ................................ . . . . 111  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   892 | 0---------    | ................................ . . . . 111  . . . .  . .. .. .. .. . .  . . . .......... ... .      |
--   893 | ----------    | ................................ . . . . ...  . . . .  . .. .. .. .. . .  . . . .......... .1. .      |
--      *=======================================================================================================================*
--
-- Table ROM32_INSTR Signal Assignments for Product Terms
MQQ962:ROM32_INSTR_PT(1) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100000000"));
MQQ963:ROM32_INSTR_PT(2) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000000"));
MQQ964:ROM32_INSTR_PT(3) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000000"));
MQQ965:ROM32_INSTR_PT(4) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000000"));
MQQ966:ROM32_INSTR_PT(5) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110000000"));
MQQ967:ROM32_INSTR_PT(6) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000000"));
MQQ968:ROM32_INSTR_PT(7) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00100000"));
MQQ969:ROM32_INSTR_PT(8) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100000"));
MQQ970:ROM32_INSTR_PT(9) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100000"));
MQQ971:ROM32_INSTR_PT(10) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100000"));
MQQ972:ROM32_INSTR_PT(11) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000000"));
MQQ973:ROM32_INSTR_PT(12) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000000"));
MQQ974:ROM32_INSTR_PT(13) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010000"));
MQQ975:ROM32_INSTR_PT(14) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010000"));
MQQ976:ROM32_INSTR_PT(15) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101010000"));
MQQ977:ROM32_INSTR_PT(16) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110000"));
MQQ978:ROM32_INSTR_PT(17) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110000"));
MQQ979:ROM32_INSTR_PT(18) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110000"));
MQQ980:ROM32_INSTR_PT(19) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110000"));
MQQ981:ROM32_INSTR_PT(20) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ982:ROM32_INSTR_PT(21) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010000"));
MQQ983:ROM32_INSTR_PT(22) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110000"));
MQQ984:ROM32_INSTR_PT(23) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ985:ROM32_INSTR_PT(24) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000000"));
MQQ986:ROM32_INSTR_PT(25) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100000"));
MQQ987:ROM32_INSTR_PT(26) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010000"));
MQQ988:ROM32_INSTR_PT(27) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010000"));
MQQ989:ROM32_INSTR_PT(28) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110000"));
MQQ990:ROM32_INSTR_PT(29) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ991:ROM32_INSTR_PT(30) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110000"));
MQQ992:ROM32_INSTR_PT(31) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010000"));
MQQ993:ROM32_INSTR_PT(32) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010000"));
MQQ994:ROM32_INSTR_PT(33) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110000"));
MQQ995:ROM32_INSTR_PT(34) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001000"));
MQQ996:ROM32_INSTR_PT(35) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001000"));
MQQ997:ROM32_INSTR_PT(36) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101001000"));
MQQ998:ROM32_INSTR_PT(37) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110001000"));
MQQ999:ROM32_INSTR_PT(38) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001000"));
MQQ1000:ROM32_INSTR_PT(39) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100101000"));
MQQ1001:ROM32_INSTR_PT(40) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101000"));
MQQ1002:ROM32_INSTR_PT(41) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001101000"));
MQQ1003:ROM32_INSTR_PT(42) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101000"));
MQQ1004:ROM32_INSTR_PT(43) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101000"));
MQQ1005:ROM32_INSTR_PT(44) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101000"));
MQQ1006:ROM32_INSTR_PT(45) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111101000"));
MQQ1007:ROM32_INSTR_PT(46) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001000"));
MQQ1008:ROM32_INSTR_PT(47) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101000"));
MQQ1009:ROM32_INSTR_PT(48) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001011000"));
MQQ1010:ROM32_INSTR_PT(49) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011011000"));
MQQ1011:ROM32_INSTR_PT(50) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011011000"));
MQQ1012:ROM32_INSTR_PT(51) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111000"));
MQQ1013:ROM32_INSTR_PT(52) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111000"));
MQQ1014:ROM32_INSTR_PT(53) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111000"));
MQQ1015:ROM32_INSTR_PT(54) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011000"));
MQQ1016:ROM32_INSTR_PT(55) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111000"));
MQQ1017:ROM32_INSTR_PT(56) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111000"));
MQQ1018:ROM32_INSTR_PT(57) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111000"));
MQQ1019:ROM32_INSTR_PT(58) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111000"));
MQQ1020:ROM32_INSTR_PT(59) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001000"));
MQQ1021:ROM32_INSTR_PT(60) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001000"));
MQQ1022:ROM32_INSTR_PT(61) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011000"));
MQQ1023:ROM32_INSTR_PT(62) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011000"));
MQQ1024:ROM32_INSTR_PT(63) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100111000"));
MQQ1025:ROM32_INSTR_PT(64) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111000"));
MQQ1026:ROM32_INSTR_PT(65) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000000"));
MQQ1027:ROM32_INSTR_PT(66) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000000"));
MQQ1028:ROM32_INSTR_PT(67) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000000"));
MQQ1029:ROM32_INSTR_PT(68) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000000"));
MQQ1030:ROM32_INSTR_PT(69) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010000"));
MQQ1031:ROM32_INSTR_PT(70) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010000"));
MQQ1032:ROM32_INSTR_PT(71) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ1033:ROM32_INSTR_PT(72) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010000"));
MQQ1034:ROM32_INSTR_PT(73) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001000"));
MQQ1035:ROM32_INSTR_PT(74) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011000"));
MQQ1036:ROM32_INSTR_PT(75) <=
    Eq(( ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000"));
MQQ1037:ROM32_INSTR_PT(76) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000100"));
MQQ1038:ROM32_INSTR_PT(77) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000100"));
MQQ1039:ROM32_INSTR_PT(78) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000100"));
MQQ1040:ROM32_INSTR_PT(79) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000100"));
MQQ1041:ROM32_INSTR_PT(80) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000100"));
MQQ1042:ROM32_INSTR_PT(81) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000100"));
MQQ1043:ROM32_INSTR_PT(82) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100100"));
MQQ1044:ROM32_INSTR_PT(83) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100100"));
MQQ1045:ROM32_INSTR_PT(84) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100100"));
MQQ1046:ROM32_INSTR_PT(85) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11100100"));
MQQ1047:ROM32_INSTR_PT(86) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100100"));
MQQ1048:ROM32_INSTR_PT(87) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000100"));
MQQ1049:ROM32_INSTR_PT(88) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000100"));
MQQ1050:ROM32_INSTR_PT(89) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100100"));
MQQ1051:ROM32_INSTR_PT(90) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110010100"));
MQQ1052:ROM32_INSTR_PT(91) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010100"));
MQQ1053:ROM32_INSTR_PT(92) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010100"));
MQQ1054:ROM32_INSTR_PT(93) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010100"));
MQQ1055:ROM32_INSTR_PT(94) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110100"));
MQQ1056:ROM32_INSTR_PT(95) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110100"));
MQQ1057:ROM32_INSTR_PT(96) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110100"));
MQQ1058:ROM32_INSTR_PT(97) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110100"));
MQQ1059:ROM32_INSTR_PT(98) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010100"));
MQQ1060:ROM32_INSTR_PT(99) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110100"));
MQQ1061:ROM32_INSTR_PT(100) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110100"));
MQQ1062:ROM32_INSTR_PT(101) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110100"));
MQQ1063:ROM32_INSTR_PT(102) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000100"));
MQQ1064:ROM32_INSTR_PT(103) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000100"));
MQQ1065:ROM32_INSTR_PT(104) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010100"));
MQQ1066:ROM32_INSTR_PT(105) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110100"));
MQQ1067:ROM32_INSTR_PT(106) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010100"));
MQQ1068:ROM32_INSTR_PT(107) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110100"));
MQQ1069:ROM32_INSTR_PT(108) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001001100"));
MQQ1070:ROM32_INSTR_PT(109) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001001100"));
MQQ1071:ROM32_INSTR_PT(110) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001100"));
MQQ1072:ROM32_INSTR_PT(111) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001100"));
MQQ1073:ROM32_INSTR_PT(112) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001100"));
MQQ1074:ROM32_INSTR_PT(113) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101100"));
MQQ1075:ROM32_INSTR_PT(114) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100101100"));
MQQ1076:ROM32_INSTR_PT(115) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010101100"));
MQQ1077:ROM32_INSTR_PT(116) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101100"));
MQQ1078:ROM32_INSTR_PT(117) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101100"));
MQQ1079:ROM32_INSTR_PT(118) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ1080:ROM32_INSTR_PT(119) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ1081:ROM32_INSTR_PT(120) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011100"));
MQQ1082:ROM32_INSTR_PT(121) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011100"));
MQQ1083:ROM32_INSTR_PT(122) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011011100"));
MQQ1084:ROM32_INSTR_PT(123) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ1085:ROM32_INSTR_PT(124) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111100"));
MQQ1086:ROM32_INSTR_PT(125) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ1087:ROM32_INSTR_PT(126) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ1088:ROM32_INSTR_PT(127) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011100"));
MQQ1089:ROM32_INSTR_PT(128) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111100"));
MQQ1090:ROM32_INSTR_PT(129) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ1091:ROM32_INSTR_PT(130) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ1092:ROM32_INSTR_PT(131) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001100"));
MQQ1093:ROM32_INSTR_PT(132) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101100"));
MQQ1094:ROM32_INSTR_PT(133) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ1095:ROM32_INSTR_PT(134) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111100"));
MQQ1096:ROM32_INSTR_PT(135) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111100"));
MQQ1097:ROM32_INSTR_PT(136) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011100"));
MQQ1098:ROM32_INSTR_PT(137) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0100100"));
MQQ1099:ROM32_INSTR_PT(138) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010100"));
MQQ1100:ROM32_INSTR_PT(139) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010100"));
MQQ1101:ROM32_INSTR_PT(140) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001100"));
MQQ1102:ROM32_INSTR_PT(141) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001100"));
MQQ1103:ROM32_INSTR_PT(142) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ1104:ROM32_INSTR_PT(143) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011100"));
MQQ1105:ROM32_INSTR_PT(144) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ1106:ROM32_INSTR_PT(145) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101100"));
MQQ1107:ROM32_INSTR_PT(146) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001100"));
MQQ1108:ROM32_INSTR_PT(147) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000000"));
MQQ1109:ROM32_INSTR_PT(148) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010000"));
MQQ1110:ROM32_INSTR_PT(149) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010000"));
MQQ1111:ROM32_INSTR_PT(150) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001000"));
MQQ1112:ROM32_INSTR_PT(151) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001000"));
MQQ1113:ROM32_INSTR_PT(152) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1000"));
MQQ1114:ROM32_INSTR_PT(153) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000100"));
MQQ1115:ROM32_INSTR_PT(154) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000100"));
MQQ1116:ROM32_INSTR_PT(155) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100100"));
MQQ1117:ROM32_INSTR_PT(156) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("00100"));
MQQ1118:ROM32_INSTR_PT(157) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010100"));
MQQ1119:ROM32_INSTR_PT(158) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ1120:ROM32_INSTR_PT(159) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ1121:ROM32_INSTR_PT(160) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011100"));
MQQ1122:ROM32_INSTR_PT(161) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111100"));
MQQ1123:ROM32_INSTR_PT(162) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011100"));
MQQ1124:ROM32_INSTR_PT(163) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111100"));
MQQ1125:ROM32_INSTR_PT(164) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000100"));
MQQ1126:ROM32_INSTR_PT(165) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101100"));
MQQ1127:ROM32_INSTR_PT(166) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ1128:ROM32_INSTR_PT(167) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("01100"));
MQQ1129:ROM32_INSTR_PT(168) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("10100"));
MQQ1130:ROM32_INSTR_PT(169) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000010"));
MQQ1131:ROM32_INSTR_PT(170) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000010"));
MQQ1132:ROM32_INSTR_PT(171) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000010"));
MQQ1133:ROM32_INSTR_PT(172) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000010"));
MQQ1134:ROM32_INSTR_PT(173) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100010"));
MQQ1135:ROM32_INSTR_PT(174) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100010"));
MQQ1136:ROM32_INSTR_PT(175) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000010"));
MQQ1137:ROM32_INSTR_PT(176) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ1138:ROM32_INSTR_PT(177) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010010"));
MQQ1139:ROM32_INSTR_PT(178) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110010"));
MQQ1140:ROM32_INSTR_PT(179) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001110010"));
MQQ1141:ROM32_INSTR_PT(180) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110010"));
MQQ1142:ROM32_INSTR_PT(181) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ1143:ROM32_INSTR_PT(182) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010010"));
MQQ1144:ROM32_INSTR_PT(183) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010010"));
MQQ1145:ROM32_INSTR_PT(184) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110010"));
MQQ1146:ROM32_INSTR_PT(185) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110010"));
MQQ1147:ROM32_INSTR_PT(186) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ1148:ROM32_INSTR_PT(187) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000010"));
MQQ1149:ROM32_INSTR_PT(188) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000010"));
MQQ1150:ROM32_INSTR_PT(189) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100010"));
MQQ1151:ROM32_INSTR_PT(190) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ1152:ROM32_INSTR_PT(191) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("000010"));
MQQ1153:ROM32_INSTR_PT(192) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010010"));
MQQ1154:ROM32_INSTR_PT(193) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110010"));
MQQ1155:ROM32_INSTR_PT(194) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110010"));
MQQ1156:ROM32_INSTR_PT(195) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110010"));
MQQ1157:ROM32_INSTR_PT(196) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ1158:ROM32_INSTR_PT(197) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110010"));
MQQ1159:ROM32_INSTR_PT(198) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ1160:ROM32_INSTR_PT(199) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001010"));
MQQ1161:ROM32_INSTR_PT(200) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001010"));
MQQ1162:ROM32_INSTR_PT(201) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101001010"));
MQQ1163:ROM32_INSTR_PT(202) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001001010"));
MQQ1164:ROM32_INSTR_PT(203) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001010"));
MQQ1165:ROM32_INSTR_PT(204) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001010"));
MQQ1166:ROM32_INSTR_PT(205) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100101010"));
MQQ1167:ROM32_INSTR_PT(206) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101010"));
MQQ1168:ROM32_INSTR_PT(207) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101010"));
MQQ1169:ROM32_INSTR_PT(208) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101010"));
MQQ1170:ROM32_INSTR_PT(209) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101010"));
MQQ1171:ROM32_INSTR_PT(210) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101010"));
MQQ1172:ROM32_INSTR_PT(211) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001010"));
MQQ1173:ROM32_INSTR_PT(212) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011010"));
MQQ1174:ROM32_INSTR_PT(213) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ1175:ROM32_INSTR_PT(214) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011010"));
MQQ1176:ROM32_INSTR_PT(215) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011011010"));
MQQ1177:ROM32_INSTR_PT(216) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111010"));
MQQ1178:ROM32_INSTR_PT(217) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111010"));
MQQ1179:ROM32_INSTR_PT(218) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011111010"));
MQQ1180:ROM32_INSTR_PT(219) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111010"));
MQQ1181:ROM32_INSTR_PT(220) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111010"));
MQQ1182:ROM32_INSTR_PT(221) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011010"));
MQQ1183:ROM32_INSTR_PT(222) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100111010"));
MQQ1184:ROM32_INSTR_PT(223) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111010"));
MQQ1185:ROM32_INSTR_PT(224) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111010"));
MQQ1186:ROM32_INSTR_PT(225) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101010"));
MQQ1187:ROM32_INSTR_PT(226) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011010"));
MQQ1188:ROM32_INSTR_PT(227) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ1189:ROM32_INSTR_PT(228) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100010"));
MQQ1190:ROM32_INSTR_PT(229) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100010"));
MQQ1191:ROM32_INSTR_PT(230) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ1192:ROM32_INSTR_PT(231) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001010"));
MQQ1193:ROM32_INSTR_PT(232) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001010"));
MQQ1194:ROM32_INSTR_PT(233) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101010"));
MQQ1195:ROM32_INSTR_PT(234) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011010"));
MQQ1196:ROM32_INSTR_PT(235) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011010"));
MQQ1197:ROM32_INSTR_PT(236) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011010"));
MQQ1198:ROM32_INSTR_PT(237) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110000110"));
MQQ1199:ROM32_INSTR_PT(238) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000110"));
MQQ1200:ROM32_INSTR_PT(239) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000110"));
MQQ1201:ROM32_INSTR_PT(240) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000110"));
MQQ1202:ROM32_INSTR_PT(241) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000110"));
MQQ1203:ROM32_INSTR_PT(242) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111000110"));
MQQ1204:ROM32_INSTR_PT(243) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000110"));
MQQ1205:ROM32_INSTR_PT(244) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000100110"));
MQQ1206:ROM32_INSTR_PT(245) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001100110"));
MQQ1207:ROM32_INSTR_PT(246) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000110"));
MQQ1208:ROM32_INSTR_PT(247) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000110"));
MQQ1209:ROM32_INSTR_PT(248) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100110"));
MQQ1210:ROM32_INSTR_PT(249) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100110"));
MQQ1211:ROM32_INSTR_PT(250) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110010110"));
MQQ1212:ROM32_INSTR_PT(251) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010110"));
MQQ1213:ROM32_INSTR_PT(252) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010110"));
MQQ1214:ROM32_INSTR_PT(253) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110110"));
MQQ1215:ROM32_INSTR_PT(254) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110110"));
MQQ1216:ROM32_INSTR_PT(255) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100110110"));
MQQ1217:ROM32_INSTR_PT(256) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110110"));
MQQ1218:ROM32_INSTR_PT(257) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110110"));
MQQ1219:ROM32_INSTR_PT(258) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100110"));
MQQ1220:ROM32_INSTR_PT(259) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010110"));
MQQ1221:ROM32_INSTR_PT(260) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100110110"));
MQQ1222:ROM32_INSTR_PT(261) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110110"));
MQQ1223:ROM32_INSTR_PT(262) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110110"));
MQQ1224:ROM32_INSTR_PT(263) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010110"));
MQQ1225:ROM32_INSTR_PT(264) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100001110"));
MQQ1226:ROM32_INSTR_PT(265) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001110"));
MQQ1227:ROM32_INSTR_PT(266) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110001110"));
MQQ1228:ROM32_INSTR_PT(267) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001110"));
MQQ1229:ROM32_INSTR_PT(268) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001110"));
MQQ1230:ROM32_INSTR_PT(269) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000101110"));
MQQ1231:ROM32_INSTR_PT(270) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100101110"));
MQQ1232:ROM32_INSTR_PT(271) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101110"));
MQQ1233:ROM32_INSTR_PT(272) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101110"));
MQQ1234:ROM32_INSTR_PT(273) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101110"));
MQQ1235:ROM32_INSTR_PT(274) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101110"));
MQQ1236:ROM32_INSTR_PT(275) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011110"));
MQQ1237:ROM32_INSTR_PT(276) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011110"));
MQQ1238:ROM32_INSTR_PT(277) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ1239:ROM32_INSTR_PT(278) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111110"));
MQQ1240:ROM32_INSTR_PT(279) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111110"));
MQQ1241:ROM32_INSTR_PT(280) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111110"));
MQQ1242:ROM32_INSTR_PT(281) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011110"));
MQQ1243:ROM32_INSTR_PT(282) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ1244:ROM32_INSTR_PT(283) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111110"));
MQQ1245:ROM32_INSTR_PT(284) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111110"));
MQQ1246:ROM32_INSTR_PT(285) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111110"));
MQQ1247:ROM32_INSTR_PT(286) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111110"));
MQQ1248:ROM32_INSTR_PT(287) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111110"));
MQQ1249:ROM32_INSTR_PT(288) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ1250:ROM32_INSTR_PT(289) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110110"));
MQQ1251:ROM32_INSTR_PT(290) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110110"));
MQQ1252:ROM32_INSTR_PT(291) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100110"));
MQQ1253:ROM32_INSTR_PT(292) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001110"));
MQQ1254:ROM32_INSTR_PT(293) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ1255:ROM32_INSTR_PT(294) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ1256:ROM32_INSTR_PT(295) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111110"));
MQQ1257:ROM32_INSTR_PT(296) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101110"));
MQQ1258:ROM32_INSTR_PT(297) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011110"));
MQQ1259:ROM32_INSTR_PT(298) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ1260:ROM32_INSTR_PT(299) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101110"));
MQQ1261:ROM32_INSTR_PT(300) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000010"));
MQQ1262:ROM32_INSTR_PT(301) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ1263:ROM32_INSTR_PT(302) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011010"));
MQQ1264:ROM32_INSTR_PT(303) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ1265:ROM32_INSTR_PT(304) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ1266:ROM32_INSTR_PT(305) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101010"));
MQQ1267:ROM32_INSTR_PT(306) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000110"));
MQQ1268:ROM32_INSTR_PT(307) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000110"));
MQQ1269:ROM32_INSTR_PT(308) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010110"));
MQQ1270:ROM32_INSTR_PT(309) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110110"));
MQQ1271:ROM32_INSTR_PT(310) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001110"));
MQQ1272:ROM32_INSTR_PT(311) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001110"));
MQQ1273:ROM32_INSTR_PT(312) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111110"));
MQQ1274:ROM32_INSTR_PT(313) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ1275:ROM32_INSTR_PT(314) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010110"));
MQQ1276:ROM32_INSTR_PT(315) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101110"));
MQQ1277:ROM32_INSTR_PT(316) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010010"));
MQQ1278:ROM32_INSTR_PT(317) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011010"));
MQQ1279:ROM32_INSTR_PT(318) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ1280:ROM32_INSTR_PT(319) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0000010"));
MQQ1281:ROM32_INSTR_PT(320) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000000"));
MQQ1282:ROM32_INSTR_PT(321) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010000"));
MQQ1283:ROM32_INSTR_PT(322) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101000"));
MQQ1284:ROM32_INSTR_PT(323) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101000"));
MQQ1285:ROM32_INSTR_PT(324) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101000"));
MQQ1286:ROM32_INSTR_PT(325) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100000"));
MQQ1287:ROM32_INSTR_PT(326) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0000100"));
MQQ1288:ROM32_INSTR_PT(327) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000100"));
MQQ1289:ROM32_INSTR_PT(328) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000100"));
MQQ1290:ROM32_INSTR_PT(329) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000100"));
MQQ1291:ROM32_INSTR_PT(330) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0100100"));
MQQ1292:ROM32_INSTR_PT(331) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001100"));
MQQ1293:ROM32_INSTR_PT(332) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00101100"));
MQQ1294:ROM32_INSTR_PT(333) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011100"));
MQQ1295:ROM32_INSTR_PT(334) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000000"));
MQQ1296:ROM32_INSTR_PT(335) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ1297:ROM32_INSTR_PT(336) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ1298:ROM32_INSTR_PT(337) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010010"));
MQQ1299:ROM32_INSTR_PT(338) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ1300:ROM32_INSTR_PT(339) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ1301:ROM32_INSTR_PT(340) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001010"));
MQQ1302:ROM32_INSTR_PT(341) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001010"));
MQQ1303:ROM32_INSTR_PT(342) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100110"));
MQQ1304:ROM32_INSTR_PT(343) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ1305:ROM32_INSTR_PT(344) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ1306:ROM32_INSTR_PT(345) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101110"));
MQQ1307:ROM32_INSTR_PT(346) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ1308:ROM32_INSTR_PT(347) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011110"));
MQQ1309:ROM32_INSTR_PT(348) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ1310:ROM32_INSTR_PT(349) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100110"));
MQQ1311:ROM32_INSTR_PT(350) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011110"));
MQQ1312:ROM32_INSTR_PT(351) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000000"));
MQQ1313:ROM32_INSTR_PT(352) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101000"));
MQQ1314:ROM32_INSTR_PT(353) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ1315:ROM32_INSTR_PT(354) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000010"));
MQQ1316:ROM32_INSTR_PT(355) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100010"));
MQQ1317:ROM32_INSTR_PT(356) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110110"));
MQQ1318:ROM32_INSTR_PT(357) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011110"));
MQQ1319:ROM32_INSTR_PT(358) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100010"));
MQQ1320:ROM32_INSTR_PT(359) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000001"));
MQQ1321:ROM32_INSTR_PT(360) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000001"));
MQQ1322:ROM32_INSTR_PT(361) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110000001"));
MQQ1323:ROM32_INSTR_PT(362) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000001"));
MQQ1324:ROM32_INSTR_PT(363) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100001"));
MQQ1325:ROM32_INSTR_PT(364) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11100001"));
MQQ1326:ROM32_INSTR_PT(365) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000001"));
MQQ1327:ROM32_INSTR_PT(366) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ1328:ROM32_INSTR_PT(367) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010001"));
MQQ1329:ROM32_INSTR_PT(368) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010001"));
MQQ1330:ROM32_INSTR_PT(369) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110001"));
MQQ1331:ROM32_INSTR_PT(370) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110001"));
MQQ1332:ROM32_INSTR_PT(371) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001110001"));
MQQ1333:ROM32_INSTR_PT(372) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00110001"));
MQQ1334:ROM32_INSTR_PT(373) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110001"));
MQQ1335:ROM32_INSTR_PT(374) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110001"));
MQQ1336:ROM32_INSTR_PT(375) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110001"));
MQQ1337:ROM32_INSTR_PT(376) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110001"));
MQQ1338:ROM32_INSTR_PT(377) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110001"));
MQQ1339:ROM32_INSTR_PT(378) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000001"));
MQQ1340:ROM32_INSTR_PT(379) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ1341:ROM32_INSTR_PT(380) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0100001"));
MQQ1342:ROM32_INSTR_PT(381) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100001"));
MQQ1343:ROM32_INSTR_PT(382) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010001"));
MQQ1344:ROM32_INSTR_PT(383) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100110001"));
MQQ1345:ROM32_INSTR_PT(384) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110001"));
MQQ1346:ROM32_INSTR_PT(385) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010001"));
MQQ1347:ROM32_INSTR_PT(386) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001001"));
MQQ1348:ROM32_INSTR_PT(387) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001001"));
MQQ1349:ROM32_INSTR_PT(388) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111001001"));
MQQ1350:ROM32_INSTR_PT(389) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001001"));
MQQ1351:ROM32_INSTR_PT(390) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001001"));
MQQ1352:ROM32_INSTR_PT(391) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101001"));
MQQ1353:ROM32_INSTR_PT(392) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100101001"));
MQQ1354:ROM32_INSTR_PT(393) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101001"));
MQQ1355:ROM32_INSTR_PT(394) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001101001"));
MQQ1356:ROM32_INSTR_PT(395) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101001"));
MQQ1357:ROM32_INSTR_PT(396) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101001"));
MQQ1358:ROM32_INSTR_PT(397) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111101001"));
MQQ1359:ROM32_INSTR_PT(398) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011001"));
MQQ1360:ROM32_INSTR_PT(399) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001011001"));
MQQ1361:ROM32_INSTR_PT(400) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011111001"));
MQQ1362:ROM32_INSTR_PT(401) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111001"));
MQQ1363:ROM32_INSTR_PT(402) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011001"));
MQQ1364:ROM32_INSTR_PT(403) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011001"));
MQQ1365:ROM32_INSTR_PT(404) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111001"));
MQQ1366:ROM32_INSTR_PT(405) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111001"));
MQQ1367:ROM32_INSTR_PT(406) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111001"));
MQQ1368:ROM32_INSTR_PT(407) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011001"));
MQQ1369:ROM32_INSTR_PT(408) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111001"));
MQQ1370:ROM32_INSTR_PT(409) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111001"));
MQQ1371:ROM32_INSTR_PT(410) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011001"));
MQQ1372:ROM32_INSTR_PT(411) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000001"));
MQQ1373:ROM32_INSTR_PT(412) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ1374:ROM32_INSTR_PT(413) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100001"));
MQQ1375:ROM32_INSTR_PT(414) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0010001"));
MQQ1376:ROM32_INSTR_PT(415) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010001"));
MQQ1377:ROM32_INSTR_PT(416) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001001"));
MQQ1378:ROM32_INSTR_PT(417) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101001"));
MQQ1379:ROM32_INSTR_PT(418) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011001"));
MQQ1380:ROM32_INSTR_PT(419) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011001"));
MQQ1381:ROM32_INSTR_PT(420) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000101"));
MQQ1382:ROM32_INSTR_PT(421) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000101"));
MQQ1383:ROM32_INSTR_PT(422) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000101"));
MQQ1384:ROM32_INSTR_PT(423) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000101"));
MQQ1385:ROM32_INSTR_PT(424) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000101"));
MQQ1386:ROM32_INSTR_PT(425) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000101"));
MQQ1387:ROM32_INSTR_PT(426) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100101"));
MQQ1388:ROM32_INSTR_PT(427) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100101"));
MQQ1389:ROM32_INSTR_PT(428) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100101"));
MQQ1390:ROM32_INSTR_PT(429) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001100101"));
MQQ1391:ROM32_INSTR_PT(430) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100101"));
MQQ1392:ROM32_INSTR_PT(431) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11100101"));
MQQ1393:ROM32_INSTR_PT(432) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100101"));
MQQ1394:ROM32_INSTR_PT(433) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110010101"));
MQQ1395:ROM32_INSTR_PT(434) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010101"));
MQQ1396:ROM32_INSTR_PT(435) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101010101"));
MQQ1397:ROM32_INSTR_PT(436) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010101"));
MQQ1398:ROM32_INSTR_PT(437) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110101"));
MQQ1399:ROM32_INSTR_PT(438) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110101"));
MQQ1400:ROM32_INSTR_PT(439) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110101"));
MQQ1401:ROM32_INSTR_PT(440) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110101"));
MQQ1402:ROM32_INSTR_PT(441) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110101"));
MQQ1403:ROM32_INSTR_PT(442) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000101"));
MQQ1404:ROM32_INSTR_PT(443) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000101"));
MQQ1405:ROM32_INSTR_PT(444) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100101"));
MQQ1406:ROM32_INSTR_PT(445) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010101"));
MQQ1407:ROM32_INSTR_PT(446) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110101"));
MQQ1408:ROM32_INSTR_PT(447) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110101"));
MQQ1409:ROM32_INSTR_PT(448) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010101"));
MQQ1410:ROM32_INSTR_PT(449) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100001101"));
MQQ1411:ROM32_INSTR_PT(450) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110001101"));
MQQ1412:ROM32_INSTR_PT(451) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001001101"));
MQQ1413:ROM32_INSTR_PT(452) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001101"));
MQQ1414:ROM32_INSTR_PT(453) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101101"));
MQQ1415:ROM32_INSTR_PT(454) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101101"));
MQQ1416:ROM32_INSTR_PT(455) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001101"));
MQQ1417:ROM32_INSTR_PT(456) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001101"));
MQQ1418:ROM32_INSTR_PT(457) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101101"));
MQQ1419:ROM32_INSTR_PT(458) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101101"));
MQQ1420:ROM32_INSTR_PT(459) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011101"));
MQQ1421:ROM32_INSTR_PT(460) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011101"));
MQQ1422:ROM32_INSTR_PT(461) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111101"));
MQQ1423:ROM32_INSTR_PT(462) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011101"));
MQQ1424:ROM32_INSTR_PT(463) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011101"));
MQQ1425:ROM32_INSTR_PT(464) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111101"));
MQQ1426:ROM32_INSTR_PT(465) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100111101"));
MQQ1427:ROM32_INSTR_PT(466) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111101"));
MQQ1428:ROM32_INSTR_PT(467) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111101"));
MQQ1429:ROM32_INSTR_PT(468) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100101"));
MQQ1430:ROM32_INSTR_PT(469) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010101"));
MQQ1431:ROM32_INSTR_PT(470) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0010101"));
MQQ1432:ROM32_INSTR_PT(471) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110101"));
MQQ1433:ROM32_INSTR_PT(472) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010101"));
MQQ1434:ROM32_INSTR_PT(473) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001101"));
MQQ1435:ROM32_INSTR_PT(474) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001101"));
MQQ1436:ROM32_INSTR_PT(475) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001101"));
MQQ1437:ROM32_INSTR_PT(476) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011101"));
MQQ1438:ROM32_INSTR_PT(477) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011101"));
MQQ1439:ROM32_INSTR_PT(478) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111101"));
MQQ1440:ROM32_INSTR_PT(479) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ1441:ROM32_INSTR_PT(480) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010001"));
MQQ1442:ROM32_INSTR_PT(481) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110001"));
MQQ1443:ROM32_INSTR_PT(482) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001001"));
MQQ1444:ROM32_INSTR_PT(483) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101001"));
MQQ1445:ROM32_INSTR_PT(484) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011001"));
MQQ1446:ROM32_INSTR_PT(485) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111001"));
MQQ1447:ROM32_INSTR_PT(486) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111001"));
MQQ1448:ROM32_INSTR_PT(487) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011001"));
MQQ1449:ROM32_INSTR_PT(488) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011001"));
MQQ1450:ROM32_INSTR_PT(489) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000101"));
MQQ1451:ROM32_INSTR_PT(490) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100101"));
MQQ1452:ROM32_INSTR_PT(491) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010101"));
MQQ1453:ROM32_INSTR_PT(492) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100101"));
MQQ1454:ROM32_INSTR_PT(493) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010101"));
MQQ1455:ROM32_INSTR_PT(494) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111101"));
MQQ1456:ROM32_INSTR_PT(495) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011101"));
MQQ1457:ROM32_INSTR_PT(496) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111101"));
MQQ1458:ROM32_INSTR_PT(497) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101101"));
MQQ1459:ROM32_INSTR_PT(498) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001101"));
MQQ1460:ROM32_INSTR_PT(499) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0000001"));
MQQ1461:ROM32_INSTR_PT(500) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001"));
MQQ1462:ROM32_INSTR_PT(501) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000011"));
MQQ1463:ROM32_INSTR_PT(502) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000011"));
MQQ1464:ROM32_INSTR_PT(503) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000011"));
MQQ1465:ROM32_INSTR_PT(504) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000011"));
MQQ1466:ROM32_INSTR_PT(505) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010100011"));
MQQ1467:ROM32_INSTR_PT(506) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100011"));
MQQ1468:ROM32_INSTR_PT(507) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100011"));
MQQ1469:ROM32_INSTR_PT(508) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000011"));
MQQ1470:ROM32_INSTR_PT(509) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100011"));
MQQ1471:ROM32_INSTR_PT(510) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000011"));
MQQ1472:ROM32_INSTR_PT(511) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010011"));
MQQ1473:ROM32_INSTR_PT(512) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010011"));
MQQ1474:ROM32_INSTR_PT(513) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010011"));
MQQ1475:ROM32_INSTR_PT(514) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010011"));
MQQ1476:ROM32_INSTR_PT(515) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010011"));
MQQ1477:ROM32_INSTR_PT(516) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101110011"));
MQQ1478:ROM32_INSTR_PT(517) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001110011"));
MQQ1479:ROM32_INSTR_PT(518) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010011"));
MQQ1480:ROM32_INSTR_PT(519) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110011"));
MQQ1481:ROM32_INSTR_PT(520) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110011"));
MQQ1482:ROM32_INSTR_PT(521) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110011"));
MQQ1483:ROM32_INSTR_PT(522) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000011"));
MQQ1484:ROM32_INSTR_PT(523) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000011"));
MQQ1485:ROM32_INSTR_PT(524) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100011"));
MQQ1486:ROM32_INSTR_PT(525) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ1487:ROM32_INSTR_PT(526) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100011"));
MQQ1488:ROM32_INSTR_PT(527) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010011"));
MQQ1489:ROM32_INSTR_PT(528) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110011"));
MQQ1490:ROM32_INSTR_PT(529) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010011"));
MQQ1491:ROM32_INSTR_PT(530) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001011"));
MQQ1492:ROM32_INSTR_PT(531) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101001011"));
MQQ1493:ROM32_INSTR_PT(532) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001001011"));
MQQ1494:ROM32_INSTR_PT(533) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111001011"));
MQQ1495:ROM32_INSTR_PT(534) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000101011"));
MQQ1496:ROM32_INSTR_PT(535) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101011"));
MQQ1497:ROM32_INSTR_PT(536) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101011"));
MQQ1498:ROM32_INSTR_PT(537) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101011"));
MQQ1499:ROM32_INSTR_PT(538) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101011"));
MQQ1500:ROM32_INSTR_PT(539) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101011"));
MQQ1501:ROM32_INSTR_PT(540) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011011"));
MQQ1502:ROM32_INSTR_PT(541) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ1503:ROM32_INSTR_PT(542) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011011"));
MQQ1504:ROM32_INSTR_PT(543) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111011"));
MQQ1505:ROM32_INSTR_PT(544) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011011"));
MQQ1506:ROM32_INSTR_PT(545) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ1507:ROM32_INSTR_PT(546) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111011"));
MQQ1508:ROM32_INSTR_PT(547) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101011"));
MQQ1509:ROM32_INSTR_PT(548) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011011"));
MQQ1510:ROM32_INSTR_PT(549) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111011"));
MQQ1511:ROM32_INSTR_PT(550) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100011"));
MQQ1512:ROM32_INSTR_PT(551) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100011"));
MQQ1513:ROM32_INSTR_PT(552) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110011"));
MQQ1514:ROM32_INSTR_PT(553) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001011"));
MQQ1515:ROM32_INSTR_PT(554) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001011"));
MQQ1516:ROM32_INSTR_PT(555) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101011"));
MQQ1517:ROM32_INSTR_PT(556) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011011"));
MQQ1518:ROM32_INSTR_PT(557) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011011"));
MQQ1519:ROM32_INSTR_PT(558) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011011"));
MQQ1520:ROM32_INSTR_PT(559) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111011"));
MQQ1521:ROM32_INSTR_PT(560) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101011"));
MQQ1522:ROM32_INSTR_PT(561) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011011"));
MQQ1523:ROM32_INSTR_PT(562) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111011"));
MQQ1524:ROM32_INSTR_PT(563) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111011"));
MQQ1525:ROM32_INSTR_PT(564) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ1526:ROM32_INSTR_PT(565) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000111"));
MQQ1527:ROM32_INSTR_PT(566) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000111"));
MQQ1528:ROM32_INSTR_PT(567) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000111"));
MQQ1529:ROM32_INSTR_PT(568) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000111"));
MQQ1530:ROM32_INSTR_PT(569) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000111"));
MQQ1531:ROM32_INSTR_PT(570) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000111"));
MQQ1532:ROM32_INSTR_PT(571) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010100111"));
MQQ1533:ROM32_INSTR_PT(572) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100111"));
MQQ1534:ROM32_INSTR_PT(573) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100111"));
MQQ1535:ROM32_INSTR_PT(574) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001100111"));
MQQ1536:ROM32_INSTR_PT(575) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100111"));
MQQ1537:ROM32_INSTR_PT(576) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000111"));
MQQ1538:ROM32_INSTR_PT(577) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000111"));
MQQ1539:ROM32_INSTR_PT(578) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010111"));
MQQ1540:ROM32_INSTR_PT(579) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010111"));
MQQ1541:ROM32_INSTR_PT(580) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001010111"));
MQQ1542:ROM32_INSTR_PT(581) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010111"));
MQQ1543:ROM32_INSTR_PT(582) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110111"));
MQQ1544:ROM32_INSTR_PT(583) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010111"));
MQQ1545:ROM32_INSTR_PT(584) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100111"));
MQQ1546:ROM32_INSTR_PT(585) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001111"));
MQQ1547:ROM32_INSTR_PT(586) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001111"));
MQQ1548:ROM32_INSTR_PT(587) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001111"));
MQQ1549:ROM32_INSTR_PT(588) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001111"));
MQQ1550:ROM32_INSTR_PT(589) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001111"));
MQQ1551:ROM32_INSTR_PT(590) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101111"));
MQQ1552:ROM32_INSTR_PT(591) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001101111"));
MQQ1553:ROM32_INSTR_PT(592) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101111"));
MQQ1554:ROM32_INSTR_PT(593) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101111"));
MQQ1555:ROM32_INSTR_PT(594) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001111"));
MQQ1556:ROM32_INSTR_PT(595) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101111"));
MQQ1557:ROM32_INSTR_PT(596) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011111"));
MQQ1558:ROM32_INSTR_PT(597) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011111"));
MQQ1559:ROM32_INSTR_PT(598) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001011111"));
MQQ1560:ROM32_INSTR_PT(599) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111111"));
MQQ1561:ROM32_INSTR_PT(600) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111111"));
MQQ1562:ROM32_INSTR_PT(601) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ1563:ROM32_INSTR_PT(602) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011111"));
MQQ1564:ROM32_INSTR_PT(603) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ1565:ROM32_INSTR_PT(604) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111111"));
MQQ1566:ROM32_INSTR_PT(605) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111111"));
MQQ1567:ROM32_INSTR_PT(606) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111111"));
MQQ1568:ROM32_INSTR_PT(607) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101111"));
MQQ1569:ROM32_INSTR_PT(608) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ1570:ROM32_INSTR_PT(609) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111111"));
MQQ1571:ROM32_INSTR_PT(610) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111111"));
MQQ1572:ROM32_INSTR_PT(611) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1573:ROM32_INSTR_PT(612) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1574:ROM32_INSTR_PT(613) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000111"));
MQQ1575:ROM32_INSTR_PT(614) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110111"));
MQQ1576:ROM32_INSTR_PT(615) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110111"));
MQQ1577:ROM32_INSTR_PT(616) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000111"));
MQQ1578:ROM32_INSTR_PT(617) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001111"));
MQQ1579:ROM32_INSTR_PT(618) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011111"));
MQQ1580:ROM32_INSTR_PT(619) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ1581:ROM32_INSTR_PT(620) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011111"));
MQQ1582:ROM32_INSTR_PT(621) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111111"));
MQQ1583:ROM32_INSTR_PT(622) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ1584:ROM32_INSTR_PT(623) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ1585:ROM32_INSTR_PT(624) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ1586:ROM32_INSTR_PT(625) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ1587:ROM32_INSTR_PT(626) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ1588:ROM32_INSTR_PT(627) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000011"));
MQQ1589:ROM32_INSTR_PT(628) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("10011"));
MQQ1590:ROM32_INSTR_PT(629) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ1591:ROM32_INSTR_PT(630) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011011"));
MQQ1592:ROM32_INSTR_PT(631) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111011"));
MQQ1593:ROM32_INSTR_PT(632) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111011"));
MQQ1594:ROM32_INSTR_PT(633) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111011"));
MQQ1595:ROM32_INSTR_PT(634) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ1596:ROM32_INSTR_PT(635) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ1597:ROM32_INSTR_PT(636) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011011"));
MQQ1598:ROM32_INSTR_PT(637) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("10011"));
MQQ1599:ROM32_INSTR_PT(638) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000111"));
MQQ1600:ROM32_INSTR_PT(639) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100111"));
MQQ1601:ROM32_INSTR_PT(640) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010111"));
MQQ1602:ROM32_INSTR_PT(641) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000111"));
MQQ1603:ROM32_INSTR_PT(642) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ1604:ROM32_INSTR_PT(643) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1605:ROM32_INSTR_PT(644) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1606:ROM32_INSTR_PT(645) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0010111"));
MQQ1607:ROM32_INSTR_PT(646) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110111"));
MQQ1608:ROM32_INSTR_PT(647) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011111"));
MQQ1609:ROM32_INSTR_PT(648) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ1610:ROM32_INSTR_PT(649) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ1611:ROM32_INSTR_PT(650) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ1612:ROM32_INSTR_PT(651) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ1613:ROM32_INSTR_PT(652) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ1614:ROM32_INSTR_PT(653) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000001"));
MQQ1615:ROM32_INSTR_PT(654) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110001"));
MQQ1616:ROM32_INSTR_PT(655) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110001"));
MQQ1617:ROM32_INSTR_PT(656) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001001"));
MQQ1618:ROM32_INSTR_PT(657) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101001"));
MQQ1619:ROM32_INSTR_PT(658) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001001"));
MQQ1620:ROM32_INSTR_PT(659) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011001"));
MQQ1621:ROM32_INSTR_PT(660) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101001"));
MQQ1622:ROM32_INSTR_PT(661) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000101"));
MQQ1623:ROM32_INSTR_PT(662) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000101"));
MQQ1624:ROM32_INSTR_PT(663) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100101"));
MQQ1625:ROM32_INSTR_PT(664) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110101"));
MQQ1626:ROM32_INSTR_PT(665) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001101"));
MQQ1627:ROM32_INSTR_PT(666) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011101"));
MQQ1628:ROM32_INSTR_PT(667) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011101"));
MQQ1629:ROM32_INSTR_PT(668) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000001"));
MQQ1630:ROM32_INSTR_PT(669) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011101"));
MQQ1631:ROM32_INSTR_PT(670) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("01001"));
MQQ1632:ROM32_INSTR_PT(671) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100101"));
MQQ1633:ROM32_INSTR_PT(672) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100011"));
MQQ1634:ROM32_INSTR_PT(673) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ1635:ROM32_INSTR_PT(674) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110011"));
MQQ1636:ROM32_INSTR_PT(675) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("000011"));
MQQ1637:ROM32_INSTR_PT(676) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ1638:ROM32_INSTR_PT(677) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101011"));
MQQ1639:ROM32_INSTR_PT(678) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011011"));
MQQ1640:ROM32_INSTR_PT(679) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011011"));
MQQ1641:ROM32_INSTR_PT(680) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ1642:ROM32_INSTR_PT(681) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010011"));
MQQ1643:ROM32_INSTR_PT(682) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100111"));
MQQ1644:ROM32_INSTR_PT(683) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010111"));
MQQ1645:ROM32_INSTR_PT(684) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010111"));
MQQ1646:ROM32_INSTR_PT(685) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001111"));
MQQ1647:ROM32_INSTR_PT(686) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101111"));
MQQ1648:ROM32_INSTR_PT(687) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011111"));
MQQ1649:ROM32_INSTR_PT(688) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ1650:ROM32_INSTR_PT(689) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ1651:ROM32_INSTR_PT(690) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1652:ROM32_INSTR_PT(691) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000111"));
MQQ1653:ROM32_INSTR_PT(692) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110111"));
MQQ1654:ROM32_INSTR_PT(693) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011111"));
MQQ1655:ROM32_INSTR_PT(694) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ1656:ROM32_INSTR_PT(695) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0011"));
MQQ1657:ROM32_INSTR_PT(696) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ1658:ROM32_INSTR_PT(697) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1659:ROM32_INSTR_PT(698) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101111"));
MQQ1660:ROM32_INSTR_PT(699) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ1661:ROM32_INSTR_PT(700) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ1662:ROM32_INSTR_PT(701) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("01111"));
MQQ1663:ROM32_INSTR_PT(702) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000001"));
MQQ1664:ROM32_INSTR_PT(703) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001001"));
MQQ1665:ROM32_INSTR_PT(704) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111001"));
MQQ1666:ROM32_INSTR_PT(705) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100001"));
MQQ1667:ROM32_INSTR_PT(706) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("001001"));
MQQ1668:ROM32_INSTR_PT(707) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111101"));
MQQ1669:ROM32_INSTR_PT(708) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0110111"));
MQQ1670:ROM32_INSTR_PT(709) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1671:ROM32_INSTR_PT(710) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ1672:ROM32_INSTR_PT(711) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1673:ROM32_INSTR_PT(712) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100111"));
MQQ1674:ROM32_INSTR_PT(713) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011111"));
MQQ1675:ROM32_INSTR_PT(714) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ1676:ROM32_INSTR_PT(715) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100101"));
MQQ1677:ROM32_INSTR_PT(716) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ1678:ROM32_INSTR_PT(717) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0111"));
MQQ1679:ROM32_INSTR_PT(718) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101"));
MQQ1680:ROM32_INSTR_PT(719) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100000"));
MQQ1681:ROM32_INSTR_PT(720) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100000"));
MQQ1682:ROM32_INSTR_PT(721) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1010000"));
MQQ1683:ROM32_INSTR_PT(722) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000110000"));
MQQ1684:ROM32_INSTR_PT(723) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ1685:ROM32_INSTR_PT(724) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100000"));
MQQ1686:ROM32_INSTR_PT(725) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111000"));
MQQ1687:ROM32_INSTR_PT(726) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0111000"));
MQQ1688:ROM32_INSTR_PT(727) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000100"));
MQQ1689:ROM32_INSTR_PT(728) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100100"));
MQQ1690:ROM32_INSTR_PT(729) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1100100"));
MQQ1691:ROM32_INSTR_PT(730) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1100100"));
MQQ1692:ROM32_INSTR_PT(731) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ1693:ROM32_INSTR_PT(732) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ1694:ROM32_INSTR_PT(733) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("10011100"));
MQQ1695:ROM32_INSTR_PT(734) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101100"));
MQQ1696:ROM32_INSTR_PT(735) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01100"));
MQQ1697:ROM32_INSTR_PT(736) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100100"));
MQQ1698:ROM32_INSTR_PT(737) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100000"));
MQQ1699:ROM32_INSTR_PT(738) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1100000"));
MQQ1700:ROM32_INSTR_PT(739) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00000100"));
MQQ1701:ROM32_INSTR_PT(740) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0101100"));
MQQ1702:ROM32_INSTR_PT(741) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011100"));
MQQ1703:ROM32_INSTR_PT(742) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ1704:ROM32_INSTR_PT(743) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11100"));
MQQ1705:ROM32_INSTR_PT(744) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000"));
MQQ1706:ROM32_INSTR_PT(745) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100010"));
MQQ1707:ROM32_INSTR_PT(746) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000010"));
MQQ1708:ROM32_INSTR_PT(747) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00010010"));
MQQ1709:ROM32_INSTR_PT(748) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00000010"));
MQQ1710:ROM32_INSTR_PT(749) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11001010"));
MQQ1711:ROM32_INSTR_PT(750) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111010"));
MQQ1712:ROM32_INSTR_PT(751) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01001010"));
MQQ1713:ROM32_INSTR_PT(752) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101010"));
MQQ1714:ROM32_INSTR_PT(753) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("010000110"));
MQQ1715:ROM32_INSTR_PT(754) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1000110"));
MQQ1716:ROM32_INSTR_PT(755) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("110100110"));
MQQ1717:ROM32_INSTR_PT(756) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0001110"));
MQQ1718:ROM32_INSTR_PT(757) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1001110"));
MQQ1719:ROM32_INSTR_PT(758) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011110"));
MQQ1720:ROM32_INSTR_PT(759) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("10011110"));
MQQ1721:ROM32_INSTR_PT(760) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ1722:ROM32_INSTR_PT(761) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("0110"));
MQQ1723:ROM32_INSTR_PT(762) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011110"));
MQQ1724:ROM32_INSTR_PT(763) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ1725:ROM32_INSTR_PT(764) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("010110"));
MQQ1726:ROM32_INSTR_PT(765) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("010100"));
MQQ1727:ROM32_INSTR_PT(766) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ1728:ROM32_INSTR_PT(767) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011100"));
MQQ1729:ROM32_INSTR_PT(768) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110000"));
MQQ1730:ROM32_INSTR_PT(769) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("00100"));
MQQ1731:ROM32_INSTR_PT(770) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100010"));
MQQ1732:ROM32_INSTR_PT(771) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1001110"));
MQQ1733:ROM32_INSTR_PT(772) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("0000"));
MQQ1734:ROM32_INSTR_PT(773) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01110"));
MQQ1735:ROM32_INSTR_PT(774) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01000001"));
MQQ1736:ROM32_INSTR_PT(775) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("110100001"));
MQQ1737:ROM32_INSTR_PT(776) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01010001"));
MQQ1738:ROM32_INSTR_PT(777) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11010001"));
MQQ1739:ROM32_INSTR_PT(778) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1010001"));
MQQ1740:ROM32_INSTR_PT(779) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000001"));
MQQ1741:ROM32_INSTR_PT(780) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1000001"));
MQQ1742:ROM32_INSTR_PT(781) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("010001"));
MQQ1743:ROM32_INSTR_PT(782) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0001001"));
MQQ1744:ROM32_INSTR_PT(783) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("001001"));
MQQ1745:ROM32_INSTR_PT(784) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011001"));
MQQ1746:ROM32_INSTR_PT(785) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111001"));
MQQ1747:ROM32_INSTR_PT(786) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011001"));
MQQ1748:ROM32_INSTR_PT(787) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00100101"));
MQQ1749:ROM32_INSTR_PT(788) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00010101"));
MQQ1750:ROM32_INSTR_PT(789) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011101"));
MQQ1751:ROM32_INSTR_PT(790) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("10011101"));
MQQ1752:ROM32_INSTR_PT(791) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011101"));
MQQ1753:ROM32_INSTR_PT(792) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110101"));
MQQ1754:ROM32_INSTR_PT(793) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("10101"));
MQQ1755:ROM32_INSTR_PT(794) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11101"));
MQQ1756:ROM32_INSTR_PT(795) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000101"));
MQQ1757:ROM32_INSTR_PT(796) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000101"));
MQQ1758:ROM32_INSTR_PT(797) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11101"));
MQQ1759:ROM32_INSTR_PT(798) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101101"));
MQQ1760:ROM32_INSTR_PT(799) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100001"));
MQQ1761:ROM32_INSTR_PT(800) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000100011"));
MQQ1762:ROM32_INSTR_PT(801) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00000011"));
MQQ1763:ROM32_INSTR_PT(802) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000011"));
MQQ1764:ROM32_INSTR_PT(803) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1010011"));
MQQ1765:ROM32_INSTR_PT(804) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("10011"));
MQQ1766:ROM32_INSTR_PT(805) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ1767:ROM32_INSTR_PT(806) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0001011"));
MQQ1768:ROM32_INSTR_PT(807) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01000011"));
MQQ1769:ROM32_INSTR_PT(808) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101011"));
MQQ1770:ROM32_INSTR_PT(809) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ1771:ROM32_INSTR_PT(810) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100111"));
MQQ1772:ROM32_INSTR_PT(811) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00010111"));
MQQ1773:ROM32_INSTR_PT(812) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01010111"));
MQQ1774:ROM32_INSTR_PT(813) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1775:ROM32_INSTR_PT(814) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1110111"));
MQQ1776:ROM32_INSTR_PT(815) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11010111"));
MQQ1777:ROM32_INSTR_PT(816) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000101111"));
MQQ1778:ROM32_INSTR_PT(817) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01101111"));
MQQ1779:ROM32_INSTR_PT(818) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1780:ROM32_INSTR_PT(819) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1781:ROM32_INSTR_PT(820) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ1782:ROM32_INSTR_PT(821) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1783:ROM32_INSTR_PT(822) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101011"));
MQQ1784:ROM32_INSTR_PT(823) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01000111"));
MQQ1785:ROM32_INSTR_PT(824) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0110111"));
MQQ1786:ROM32_INSTR_PT(825) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1787:ROM32_INSTR_PT(826) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101111"));
MQQ1788:ROM32_INSTR_PT(827) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ1789:ROM32_INSTR_PT(828) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("0111"));
MQQ1790:ROM32_INSTR_PT(829) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1791:ROM32_INSTR_PT(830) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01111"));
MQQ1792:ROM32_INSTR_PT(831) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110001"));
MQQ1793:ROM32_INSTR_PT(832) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011001"));
MQQ1794:ROM32_INSTR_PT(833) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1001101"));
MQQ1795:ROM32_INSTR_PT(834) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01001"));
MQQ1796:ROM32_INSTR_PT(835) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100011"));
MQQ1797:ROM32_INSTR_PT(836) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1111011"));
MQQ1798:ROM32_INSTR_PT(837) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ1799:ROM32_INSTR_PT(838) <=
    Eq(( ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("011"));
MQQ1800:ROM32_INSTR_PT(839) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000111"));
MQQ1801:ROM32_INSTR_PT(840) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ1802:ROM32_INSTR_PT(841) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011111"));
MQQ1803:ROM32_INSTR_PT(842) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101111"));
MQQ1804:ROM32_INSTR_PT(843) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ1805:ROM32_INSTR_PT(844) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1806:ROM32_INSTR_PT(845) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011111"));
MQQ1807:ROM32_INSTR_PT(846) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("000101"));
MQQ1808:ROM32_INSTR_PT(847) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ1809:ROM32_INSTR_PT(848) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("1111"));
MQQ1810:ROM32_INSTR_PT(849) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("10111"));
MQQ1811:ROM32_INSTR_PT(850) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("0111"));
MQQ1812:ROM32_INSTR_PT(851) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1001000"));
MQQ1813:ROM32_INSTR_PT(852) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("110000"));
MQQ1814:ROM32_INSTR_PT(853) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("00011100"));
MQQ1815:ROM32_INSTR_PT(854) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("00000010"));
MQQ1816:ROM32_INSTR_PT(855) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0100010"));
MQQ1817:ROM32_INSTR_PT(856) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0000010"));
MQQ1818:ROM32_INSTR_PT(857) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("101110"));
MQQ1819:ROM32_INSTR_PT(858) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1101110"));
MQQ1820:ROM32_INSTR_PT(859) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1001100"));
MQQ1821:ROM32_INSTR_PT(860) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("00000"));
MQQ1822:ROM32_INSTR_PT(861) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("1110"));
MQQ1823:ROM32_INSTR_PT(862) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0100101"));
MQQ1824:ROM32_INSTR_PT(863) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1001101"));
MQQ1825:ROM32_INSTR_PT(864) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("001101"));
MQQ1826:ROM32_INSTR_PT(865) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1101101"));
MQQ1827:ROM32_INSTR_PT(866) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("1101"));
MQQ1828:ROM32_INSTR_PT(867) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1010011"));
MQQ1829:ROM32_INSTR_PT(868) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1001011"));
MQQ1830:ROM32_INSTR_PT(869) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1831:ROM32_INSTR_PT(870) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0011111"));
MQQ1832:ROM32_INSTR_PT(871) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1833:ROM32_INSTR_PT(872) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1834:ROM32_INSTR_PT(873) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ1835:ROM32_INSTR_PT(874) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("01111"));
MQQ1836:ROM32_INSTR_PT(875) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("1101"));
MQQ1837:ROM32_INSTR_PT(876) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("000011"));
MQQ1838:ROM32_INSTR_PT(877) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) ) , STD_ULOGIC_VECTOR'("0000100"));
MQQ1839:ROM32_INSTR_PT(878) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6)
     ) , STD_ULOGIC_VECTOR'("010010"));
MQQ1840:ROM32_INSTR_PT(879) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(6)
     ) , STD_ULOGIC_VECTOR'("00"));
MQQ1841:ROM32_INSTR_PT(880) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) ) , STD_ULOGIC_VECTOR'("111"));
MQQ1842:ROM32_INSTR_PT(881) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1843:ROM32_INSTR_PT(882) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5)
     ) , STD_ULOGIC_VECTOR'("00"));
MQQ1844:ROM32_INSTR_PT(883) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(5)
     ) , STD_ULOGIC_VECTOR'("00"));
MQQ1845:ROM32_INSTR_PT(884) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5)
     ) , STD_ULOGIC_VECTOR'("0110"));
MQQ1846:ROM32_INSTR_PT(885) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5)
     ) , STD_ULOGIC_VECTOR'("0110"));
MQQ1847:ROM32_INSTR_PT(886) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) ) , STD_ULOGIC_VECTOR'("111"));
MQQ1848:ROM32_INSTR_PT(887) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) ) , STD_ULOGIC_VECTOR'("000"));
MQQ1849:ROM32_INSTR_PT(888) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4)
     ) , STD_ULOGIC_VECTOR'("0111"));
MQQ1850:ROM32_INSTR_PT(889) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) ) , STD_ULOGIC_VECTOR'("111"));
MQQ1851:ROM32_INSTR_PT(890) <=
    Eq(( ROM_ADDR_L2(2) ) , STD_ULOGIC'('1'));
MQQ1852:ROM32_INSTR_PT(891) <=
    Eq(( ROM_ADDR_L2(1) ) , STD_ULOGIC'('1'));
MQQ1853:ROM32_INSTR_PT(892) <=
    Eq(( ROM_ADDR_L2(0) ) , STD_ULOGIC'('0'));
MQQ1854:ROM32_INSTR_PT(893) <=
    '1';
-- Table ROM32_INSTR Signal Assignments for Outputs
MQQ1855:TEMPLATE(0) <= 
    (ROM32_INSTR_PT(28) OR ROM32_INSTR_PT(33)
     OR ROM32_INSTR_PT(45) OR ROM32_INSTR_PT(68)
     OR ROM32_INSTR_PT(76) OR ROM32_INSTR_PT(85)
     OR ROM32_INSTR_PT(113) OR ROM32_INSTR_PT(120)
     OR ROM32_INSTR_PT(128) OR ROM32_INSTR_PT(132)
     OR ROM32_INSTR_PT(142) OR ROM32_INSTR_PT(159)
     OR ROM32_INSTR_PT(162) OR ROM32_INSTR_PT(175)
     OR ROM32_INSTR_PT(176) OR ROM32_INSTR_PT(177)
     OR ROM32_INSTR_PT(180) OR ROM32_INSTR_PT(222)
     OR ROM32_INSTR_PT(226) OR ROM32_INSTR_PT(233)
     OR ROM32_INSTR_PT(237) OR ROM32_INSTR_PT(242)
     OR ROM32_INSTR_PT(255) OR ROM32_INSTR_PT(290)
     OR ROM32_INSTR_PT(292) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(335) OR ROM32_INSTR_PT(346)
     OR ROM32_INSTR_PT(351) OR ROM32_INSTR_PT(353)
     OR ROM32_INSTR_PT(356) OR ROM32_INSTR_PT(357)
     OR ROM32_INSTR_PT(359) OR ROM32_INSTR_PT(364)
     OR ROM32_INSTR_PT(365) OR ROM32_INSTR_PT(373)
     OR ROM32_INSTR_PT(381) OR ROM32_INSTR_PT(388)
     OR ROM32_INSTR_PT(391) OR ROM32_INSTR_PT(399)
     OR ROM32_INSTR_PT(425) OR ROM32_INSTR_PT(431)
     OR ROM32_INSTR_PT(467) OR ROM32_INSTR_PT(473)
     OR ROM32_INSTR_PT(527) OR ROM32_INSTR_PT(555)
     OR ROM32_INSTR_PT(563) OR ROM32_INSTR_PT(571)
     OR ROM32_INSTR_PT(586) OR ROM32_INSTR_PT(597)
     OR ROM32_INSTR_PT(604) OR ROM32_INSTR_PT(615)
     OR ROM32_INSTR_PT(652) OR ROM32_INSTR_PT(657)
     OR ROM32_INSTR_PT(664) OR ROM32_INSTR_PT(691)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(697)
     OR ROM32_INSTR_PT(711) OR ROM32_INSTR_PT(715)
     OR ROM32_INSTR_PT(716) OR ROM32_INSTR_PT(718)
     OR ROM32_INSTR_PT(729) OR ROM32_INSTR_PT(763)
     OR ROM32_INSTR_PT(792) OR ROM32_INSTR_PT(829)
     OR ROM32_INSTR_PT(831) OR ROM32_INSTR_PT(857)
     OR ROM32_INSTR_PT(872));
MQQ1856:TEMPLATE(1) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(7)
     OR ROM32_INSTR_PT(8) OR ROM32_INSTR_PT(9)
     OR ROM32_INSTR_PT(10) OR ROM32_INSTR_PT(13)
     OR ROM32_INSTR_PT(14) OR ROM32_INSTR_PT(16)
     OR ROM32_INSTR_PT(17) OR ROM32_INSTR_PT(20)
     OR ROM32_INSTR_PT(23) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(32) OR ROM32_INSTR_PT(35)
     OR ROM32_INSTR_PT(37) OR ROM32_INSTR_PT(39)
     OR ROM32_INSTR_PT(41) OR ROM32_INSTR_PT(42)
     OR ROM32_INSTR_PT(43) OR ROM32_INSTR_PT(49)
     OR ROM32_INSTR_PT(50) OR ROM32_INSTR_PT(51)
     OR ROM32_INSTR_PT(52) OR ROM32_INSTR_PT(53)
     OR ROM32_INSTR_PT(55) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(59)
     OR ROM32_INSTR_PT(63) OR ROM32_INSTR_PT(66)
     OR ROM32_INSTR_PT(67) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(73) OR ROM32_INSTR_PT(74)
     OR ROM32_INSTR_PT(77) OR ROM32_INSTR_PT(79)
     OR ROM32_INSTR_PT(80) OR ROM32_INSTR_PT(83)
     OR ROM32_INSTR_PT(84) OR ROM32_INSTR_PT(87)
     OR ROM32_INSTR_PT(90) OR ROM32_INSTR_PT(92)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(96)
     OR ROM32_INSTR_PT(97) OR ROM32_INSTR_PT(99)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(102) OR ROM32_INSTR_PT(103)
     OR ROM32_INSTR_PT(105) OR ROM32_INSTR_PT(106)
     OR ROM32_INSTR_PT(109) OR ROM32_INSTR_PT(110)
     OR ROM32_INSTR_PT(111) OR ROM32_INSTR_PT(114)
     OR ROM32_INSTR_PT(115) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(122) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(127) OR ROM32_INSTR_PT(130)
     OR ROM32_INSTR_PT(134) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(139) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(144) OR ROM32_INSTR_PT(148)
     OR ROM32_INSTR_PT(153) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(163) OR ROM32_INSTR_PT(164)
     OR ROM32_INSTR_PT(165) OR ROM32_INSTR_PT(169)
     OR ROM32_INSTR_PT(170) OR ROM32_INSTR_PT(171)
     OR ROM32_INSTR_PT(172) OR ROM32_INSTR_PT(179)
     OR ROM32_INSTR_PT(183) OR ROM32_INSTR_PT(184)
     OR ROM32_INSTR_PT(186) OR ROM32_INSTR_PT(192)
     OR ROM32_INSTR_PT(193) OR ROM32_INSTR_PT(195)
     OR ROM32_INSTR_PT(196) OR ROM32_INSTR_PT(199)
     OR ROM32_INSTR_PT(200) OR ROM32_INSTR_PT(202)
     OR ROM32_INSTR_PT(203) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(206) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(209) OR ROM32_INSTR_PT(215)
     OR ROM32_INSTR_PT(216) OR ROM32_INSTR_PT(218)
     OR ROM32_INSTR_PT(219) OR ROM32_INSTR_PT(220)
     OR ROM32_INSTR_PT(223) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(241)
     OR ROM32_INSTR_PT(243) OR ROM32_INSTR_PT(249)
     OR ROM32_INSTR_PT(250) OR ROM32_INSTR_PT(252)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(259)
     OR ROM32_INSTR_PT(260) OR ROM32_INSTR_PT(261)
     OR ROM32_INSTR_PT(262) OR ROM32_INSTR_PT(264)
     OR ROM32_INSTR_PT(267) OR ROM32_INSTR_PT(268)
     OR ROM32_INSTR_PT(269) OR ROM32_INSTR_PT(270)
     OR ROM32_INSTR_PT(273) OR ROM32_INSTR_PT(274)
     OR ROM32_INSTR_PT(275) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(280) OR ROM32_INSTR_PT(282)
     OR ROM32_INSTR_PT(283) OR ROM32_INSTR_PT(284)
     OR ROM32_INSTR_PT(287) OR ROM32_INSTR_PT(288)
     OR ROM32_INSTR_PT(289) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(306) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(321) OR ROM32_INSTR_PT(323)
     OR ROM32_INSTR_PT(328) OR ROM32_INSTR_PT(331)
     OR ROM32_INSTR_PT(342) OR ROM32_INSTR_PT(345)
     OR ROM32_INSTR_PT(348) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(352) OR ROM32_INSTR_PT(355)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(362)
     OR ROM32_INSTR_PT(363) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(368)
     OR ROM32_INSTR_PT(370) OR ROM32_INSTR_PT(371)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(382)
     OR ROM32_INSTR_PT(383) OR ROM32_INSTR_PT(386)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(390)
     OR ROM32_INSTR_PT(392) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(396) OR ROM32_INSTR_PT(400)
     OR ROM32_INSTR_PT(401) OR ROM32_INSTR_PT(402)
     OR ROM32_INSTR_PT(404) OR ROM32_INSTR_PT(405)
     OR ROM32_INSTR_PT(406) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(411) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(417)
     OR ROM32_INSTR_PT(418) OR ROM32_INSTR_PT(421)
     OR ROM32_INSTR_PT(422) OR ROM32_INSTR_PT(423)
     OR ROM32_INSTR_PT(424) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(428) OR ROM32_INSTR_PT(430)
     OR ROM32_INSTR_PT(433) OR ROM32_INSTR_PT(434)
     OR ROM32_INSTR_PT(435) OR ROM32_INSTR_PT(436)
     OR ROM32_INSTR_PT(438) OR ROM32_INSTR_PT(441)
     OR ROM32_INSTR_PT(442) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(452)
     OR ROM32_INSTR_PT(453) OR ROM32_INSTR_PT(454)
     OR ROM32_INSTR_PT(458) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(464) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(474)
     OR ROM32_INSTR_PT(475) OR ROM32_INSTR_PT(476)
     OR ROM32_INSTR_PT(477) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(480)
     OR ROM32_INSTR_PT(481) OR ROM32_INSTR_PT(482)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(491) OR ROM32_INSTR_PT(494)
     OR ROM32_INSTR_PT(496) OR ROM32_INSTR_PT(497)
     OR ROM32_INSTR_PT(498) OR ROM32_INSTR_PT(501)
     OR ROM32_INSTR_PT(502) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(505) OR ROM32_INSTR_PT(506)
     OR ROM32_INSTR_PT(507) OR ROM32_INSTR_PT(508)
     OR ROM32_INSTR_PT(509) OR ROM32_INSTR_PT(514)
     OR ROM32_INSTR_PT(517) OR ROM32_INSTR_PT(519)
     OR ROM32_INSTR_PT(520) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(524)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(531)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(535) OR ROM32_INSTR_PT(536)
     OR ROM32_INSTR_PT(538) OR ROM32_INSTR_PT(539)
     OR ROM32_INSTR_PT(541) OR ROM32_INSTR_PT(543)
     OR ROM32_INSTR_PT(544) OR ROM32_INSTR_PT(546)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(550)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(556)
     OR ROM32_INSTR_PT(557) OR ROM32_INSTR_PT(558)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(566)
     OR ROM32_INSTR_PT(568) OR ROM32_INSTR_PT(569)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(575) OR ROM32_INSTR_PT(578)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(580)
     OR ROM32_INSTR_PT(581) OR ROM32_INSTR_PT(582)
     OR ROM32_INSTR_PT(583) OR ROM32_INSTR_PT(584)
     OR ROM32_INSTR_PT(585) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(589) OR ROM32_INSTR_PT(590)
     OR ROM32_INSTR_PT(593) OR ROM32_INSTR_PT(595)
     OR ROM32_INSTR_PT(598) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(601)
     OR ROM32_INSTR_PT(602) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(606) OR ROM32_INSTR_PT(607)
     OR ROM32_INSTR_PT(608) OR ROM32_INSTR_PT(609)
     OR ROM32_INSTR_PT(610) OR ROM32_INSTR_PT(611)
     OR ROM32_INSTR_PT(612) OR ROM32_INSTR_PT(613)
     OR ROM32_INSTR_PT(614) OR ROM32_INSTR_PT(620)
     OR ROM32_INSTR_PT(621) OR ROM32_INSTR_PT(624)
     OR ROM32_INSTR_PT(625) OR ROM32_INSTR_PT(626)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(634)
     OR ROM32_INSTR_PT(635) OR ROM32_INSTR_PT(638)
     OR ROM32_INSTR_PT(639) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(643) OR ROM32_INSTR_PT(644)
     OR ROM32_INSTR_PT(647) OR ROM32_INSTR_PT(654)
     OR ROM32_INSTR_PT(660) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(666) OR ROM32_INSTR_PT(674)
     OR ROM32_INSTR_PT(677) OR ROM32_INSTR_PT(678)
     OR ROM32_INSTR_PT(680) OR ROM32_INSTR_PT(684)
     OR ROM32_INSTR_PT(685) OR ROM32_INSTR_PT(698)
     OR ROM32_INSTR_PT(708) OR ROM32_INSTR_PT(713)
     OR ROM32_INSTR_PT(719) OR ROM32_INSTR_PT(726)
     OR ROM32_INSTR_PT(733) OR ROM32_INSTR_PT(736)
     OR ROM32_INSTR_PT(745) OR ROM32_INSTR_PT(755)
     OR ROM32_INSTR_PT(762) OR ROM32_INSTR_PT(770)
     OR ROM32_INSTR_PT(785) OR ROM32_INSTR_PT(795)
     OR ROM32_INSTR_PT(801) OR ROM32_INSTR_PT(805)
     OR ROM32_INSTR_PT(812) OR ROM32_INSTR_PT(817)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(845)
     OR ROM32_INSTR_PT(847) OR ROM32_INSTR_PT(851)
     OR ROM32_INSTR_PT(853) OR ROM32_INSTR_PT(854)
     OR ROM32_INSTR_PT(855) OR ROM32_INSTR_PT(862)
     OR ROM32_INSTR_PT(869) OR ROM32_INSTR_PT(870)
     OR ROM32_INSTR_PT(871) OR ROM32_INSTR_PT(878)
     OR ROM32_INSTR_PT(889));
MQQ1857:TEMPLATE(2) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(7)
     OR ROM32_INSTR_PT(13) OR ROM32_INSTR_PT(14)
     OR ROM32_INSTR_PT(18) OR ROM32_INSTR_PT(23)
     OR ROM32_INSTR_PT(27) OR ROM32_INSTR_PT(29)
     OR ROM32_INSTR_PT(31) OR ROM32_INSTR_PT(35)
     OR ROM32_INSTR_PT(38) OR ROM32_INSTR_PT(39)
     OR ROM32_INSTR_PT(41) OR ROM32_INSTR_PT(42)
     OR ROM32_INSTR_PT(43) OR ROM32_INSTR_PT(53)
     OR ROM32_INSTR_PT(56) OR ROM32_INSTR_PT(57)
     OR ROM32_INSTR_PT(62) OR ROM32_INSTR_PT(70)
     OR ROM32_INSTR_PT(72) OR ROM32_INSTR_PT(79)
     OR ROM32_INSTR_PT(80) OR ROM32_INSTR_PT(81)
     OR ROM32_INSTR_PT(83) OR ROM32_INSTR_PT(92)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(98) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(102) OR ROM32_INSTR_PT(105)
     OR ROM32_INSTR_PT(109) OR ROM32_INSTR_PT(110)
     OR ROM32_INSTR_PT(111) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(122) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(130) OR ROM32_INSTR_PT(139)
     OR ROM32_INSTR_PT(141) OR ROM32_INSTR_PT(144)
     OR ROM32_INSTR_PT(145) OR ROM32_INSTR_PT(146)
     OR ROM32_INSTR_PT(147) OR ROM32_INSTR_PT(150)
     OR ROM32_INSTR_PT(151) OR ROM32_INSTR_PT(153)
     OR ROM32_INSTR_PT(158) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(165) OR ROM32_INSTR_PT(166)
     OR ROM32_INSTR_PT(172) OR ROM32_INSTR_PT(174)
     OR ROM32_INSTR_PT(185) OR ROM32_INSTR_PT(186)
     OR ROM32_INSTR_PT(187) OR ROM32_INSTR_PT(189)
     OR ROM32_INSTR_PT(192) OR ROM32_INSTR_PT(193)
     OR ROM32_INSTR_PT(195) OR ROM32_INSTR_PT(199)
     OR ROM32_INSTR_PT(203) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(206) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(208) OR ROM32_INSTR_PT(209)
     OR ROM32_INSTR_PT(210) OR ROM32_INSTR_PT(218)
     OR ROM32_INSTR_PT(228) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(230) OR ROM32_INSTR_PT(232)
     OR ROM32_INSTR_PT(235) OR ROM32_INSTR_PT(240)
     OR ROM32_INSTR_PT(245) OR ROM32_INSTR_PT(249)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(252)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(262)
     OR ROM32_INSTR_PT(268) OR ROM32_INSTR_PT(275)
     OR ROM32_INSTR_PT(279) OR ROM32_INSTR_PT(285)
     OR ROM32_INSTR_PT(287) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(291) OR ROM32_INSTR_PT(294)
     OR ROM32_INSTR_PT(302) OR ROM32_INSTR_PT(305)
     OR ROM32_INSTR_PT(307) OR ROM32_INSTR_PT(311)
     OR ROM32_INSTR_PT(322) OR ROM32_INSTR_PT(323)
     OR ROM32_INSTR_PT(325) OR ROM32_INSTR_PT(329)
     OR ROM32_INSTR_PT(331) OR ROM32_INSTR_PT(332)
     OR ROM32_INSTR_PT(337) OR ROM32_INSTR_PT(338)
     OR ROM32_INSTR_PT(339) OR ROM32_INSTR_PT(342)
     OR ROM32_INSTR_PT(350) OR ROM32_INSTR_PT(352)
     OR ROM32_INSTR_PT(355) OR ROM32_INSTR_PT(362)
     OR ROM32_INSTR_PT(363) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(368)
     OR ROM32_INSTR_PT(370) OR ROM32_INSTR_PT(374)
     OR ROM32_INSTR_PT(376) OR ROM32_INSTR_PT(378)
     OR ROM32_INSTR_PT(382) OR ROM32_INSTR_PT(386)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(393)
     OR ROM32_INSTR_PT(394) OR ROM32_INSTR_PT(395)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(400)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(404)
     OR ROM32_INSTR_PT(405) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(416)
     OR ROM32_INSTR_PT(417) OR ROM32_INSTR_PT(418)
     OR ROM32_INSTR_PT(419) OR ROM32_INSTR_PT(422)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(435)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(438)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(442)
     OR ROM32_INSTR_PT(443) OR ROM32_INSTR_PT(446)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(452)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(456)
     OR ROM32_INSTR_PT(458) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(463) OR ROM32_INSTR_PT(464)
     OR ROM32_INSTR_PT(465) OR ROM32_INSTR_PT(468)
     OR ROM32_INSTR_PT(469) OR ROM32_INSTR_PT(471)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(474)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(480)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(489)
     OR ROM32_INSTR_PT(496) OR ROM32_INSTR_PT(497)
     OR ROM32_INSTR_PT(498) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(505) OR ROM32_INSTR_PT(507)
     OR ROM32_INSTR_PT(513) OR ROM32_INSTR_PT(514)
     OR ROM32_INSTR_PT(517) OR ROM32_INSTR_PT(532)
     OR ROM32_INSTR_PT(537) OR ROM32_INSTR_PT(539)
     OR ROM32_INSTR_PT(541) OR ROM32_INSTR_PT(544)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(549)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(561)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(569)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(577) OR ROM32_INSTR_PT(579)
     OR ROM32_INSTR_PT(580) OR ROM32_INSTR_PT(584)
     OR ROM32_INSTR_PT(587) OR ROM32_INSTR_PT(589)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(593)
     OR ROM32_INSTR_PT(596) OR ROM32_INSTR_PT(598)
     OR ROM32_INSTR_PT(599) OR ROM32_INSTR_PT(600)
     OR ROM32_INSTR_PT(605) OR ROM32_INSTR_PT(606)
     OR ROM32_INSTR_PT(607) OR ROM32_INSTR_PT(608)
     OR ROM32_INSTR_PT(609) OR ROM32_INSTR_PT(610)
     OR ROM32_INSTR_PT(611) OR ROM32_INSTR_PT(614)
     OR ROM32_INSTR_PT(620) OR ROM32_INSTR_PT(624)
     OR ROM32_INSTR_PT(625) OR ROM32_INSTR_PT(629)
     OR ROM32_INSTR_PT(632) OR ROM32_INSTR_PT(634)
     OR ROM32_INSTR_PT(638) OR ROM32_INSTR_PT(640)
     OR ROM32_INSTR_PT(643) OR ROM32_INSTR_PT(653)
     OR ROM32_INSTR_PT(659) OR ROM32_INSTR_PT(660)
     OR ROM32_INSTR_PT(663) OR ROM32_INSTR_PT(668)
     OR ROM32_INSTR_PT(672) OR ROM32_INSTR_PT(678)
     OR ROM32_INSTR_PT(680) OR ROM32_INSTR_PT(684)
     OR ROM32_INSTR_PT(685) OR ROM32_INSTR_PT(689)
     OR ROM32_INSTR_PT(698) OR ROM32_INSTR_PT(704)
     OR ROM32_INSTR_PT(705) OR ROM32_INSTR_PT(708)
     OR ROM32_INSTR_PT(713) OR ROM32_INSTR_PT(720)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(733)
     OR ROM32_INSTR_PT(751) OR ROM32_INSTR_PT(752)
     OR ROM32_INSTR_PT(753) OR ROM32_INSTR_PT(759)
     OR ROM32_INSTR_PT(774) OR ROM32_INSTR_PT(785)
     OR ROM32_INSTR_PT(787) OR ROM32_INSTR_PT(790)
     OR ROM32_INSTR_PT(795) OR ROM32_INSTR_PT(799)
     OR ROM32_INSTR_PT(801) OR ROM32_INSTR_PT(803)
     OR ROM32_INSTR_PT(805) OR ROM32_INSTR_PT(807)
     OR ROM32_INSTR_PT(812) OR ROM32_INSTR_PT(817)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(823)
     OR ROM32_INSTR_PT(845) OR ROM32_INSTR_PT(847)
     OR ROM32_INSTR_PT(851) OR ROM32_INSTR_PT(853)
     OR ROM32_INSTR_PT(854) OR ROM32_INSTR_PT(869)
     OR ROM32_INSTR_PT(871) OR ROM32_INSTR_PT(878)
     OR ROM32_INSTR_PT(881) OR ROM32_INSTR_PT(889)
    );
MQQ1858:TEMPLATE(3) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(7)
     OR ROM32_INSTR_PT(8) OR ROM32_INSTR_PT(9)
     OR ROM32_INSTR_PT(10) OR ROM32_INSTR_PT(13)
     OR ROM32_INSTR_PT(14) OR ROM32_INSTR_PT(16)
     OR ROM32_INSTR_PT(17) OR ROM32_INSTR_PT(18)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(23)
     OR ROM32_INSTR_PT(26) OR ROM32_INSTR_PT(27)
     OR ROM32_INSTR_PT(28) OR ROM32_INSTR_PT(31)
     OR ROM32_INSTR_PT(32) OR ROM32_INSTR_PT(33)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(37)
     OR ROM32_INSTR_PT(38) OR ROM32_INSTR_PT(39)
     OR ROM32_INSTR_PT(41) OR ROM32_INSTR_PT(42)
     OR ROM32_INSTR_PT(43) OR ROM32_INSTR_PT(45)
     OR ROM32_INSTR_PT(49) OR ROM32_INSTR_PT(52)
     OR ROM32_INSTR_PT(53) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(59)
     OR ROM32_INSTR_PT(62) OR ROM32_INSTR_PT(63)
     OR ROM32_INSTR_PT(66) OR ROM32_INSTR_PT(67)
     OR ROM32_INSTR_PT(70) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(73) OR ROM32_INSTR_PT(74)
     OR ROM32_INSTR_PT(77) OR ROM32_INSTR_PT(78)
     OR ROM32_INSTR_PT(79) OR ROM32_INSTR_PT(80)
     OR ROM32_INSTR_PT(83) OR ROM32_INSTR_PT(84)
     OR ROM32_INSTR_PT(85) OR ROM32_INSTR_PT(87)
     OR ROM32_INSTR_PT(90) OR ROM32_INSTR_PT(92)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(97) OR ROM32_INSTR_PT(98)
     OR ROM32_INSTR_PT(99) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(102) OR ROM32_INSTR_PT(103)
     OR ROM32_INSTR_PT(105) OR ROM32_INSTR_PT(109)
     OR ROM32_INSTR_PT(110) OR ROM32_INSTR_PT(111)
     OR ROM32_INSTR_PT(114) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(122) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(127) OR ROM32_INSTR_PT(130)
     OR ROM32_INSTR_PT(131) OR ROM32_INSTR_PT(134)
     OR ROM32_INSTR_PT(139) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(144) OR ROM32_INSTR_PT(145)
     OR ROM32_INSTR_PT(146) OR ROM32_INSTR_PT(147)
     OR ROM32_INSTR_PT(148) OR ROM32_INSTR_PT(150)
     OR ROM32_INSTR_PT(151) OR ROM32_INSTR_PT(153)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(162) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(164) OR ROM32_INSTR_PT(165)
     OR ROM32_INSTR_PT(166) OR ROM32_INSTR_PT(169)
     OR ROM32_INSTR_PT(171) OR ROM32_INSTR_PT(172)
     OR ROM32_INSTR_PT(173) OR ROM32_INSTR_PT(174)
     OR ROM32_INSTR_PT(176) OR ROM32_INSTR_PT(177)
     OR ROM32_INSTR_PT(178) OR ROM32_INSTR_PT(179)
     OR ROM32_INSTR_PT(180) OR ROM32_INSTR_PT(181)
     OR ROM32_INSTR_PT(184) OR ROM32_INSTR_PT(185)
     OR ROM32_INSTR_PT(186) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(189) OR ROM32_INSTR_PT(192)
     OR ROM32_INSTR_PT(194) OR ROM32_INSTR_PT(199)
     OR ROM32_INSTR_PT(200) OR ROM32_INSTR_PT(202)
     OR ROM32_INSTR_PT(203) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(206) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(208) OR ROM32_INSTR_PT(209)
     OR ROM32_INSTR_PT(210) OR ROM32_INSTR_PT(212)
     OR ROM32_INSTR_PT(216) OR ROM32_INSTR_PT(218)
     OR ROM32_INSTR_PT(219) OR ROM32_INSTR_PT(220)
     OR ROM32_INSTR_PT(222) OR ROM32_INSTR_PT(223)
     OR ROM32_INSTR_PT(224) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(228)
     OR ROM32_INSTR_PT(229) OR ROM32_INSTR_PT(230)
     OR ROM32_INSTR_PT(232) OR ROM32_INSTR_PT(233)
     OR ROM32_INSTR_PT(235) OR ROM32_INSTR_PT(238)
     OR ROM32_INSTR_PT(240) OR ROM32_INSTR_PT(242)
     OR ROM32_INSTR_PT(244) OR ROM32_INSTR_PT(245)
     OR ROM32_INSTR_PT(249) OR ROM32_INSTR_PT(250)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(252)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(255)
     OR ROM32_INSTR_PT(256) OR ROM32_INSTR_PT(257)
     OR ROM32_INSTR_PT(259) OR ROM32_INSTR_PT(261)
     OR ROM32_INSTR_PT(262) OR ROM32_INSTR_PT(264)
     OR ROM32_INSTR_PT(266) OR ROM32_INSTR_PT(267)
     OR ROM32_INSTR_PT(268) OR ROM32_INSTR_PT(269)
     OR ROM32_INSTR_PT(270) OR ROM32_INSTR_PT(271)
     OR ROM32_INSTR_PT(272) OR ROM32_INSTR_PT(273)
     OR ROM32_INSTR_PT(275) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(279) OR ROM32_INSTR_PT(280)
     OR ROM32_INSTR_PT(284) OR ROM32_INSTR_PT(285)
     OR ROM32_INSTR_PT(288) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(290) OR ROM32_INSTR_PT(291)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(302)
     OR ROM32_INSTR_PT(303) OR ROM32_INSTR_PT(305)
     OR ROM32_INSTR_PT(307) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(311) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(322)
     OR ROM32_INSTR_PT(323) OR ROM32_INSTR_PT(325)
     OR ROM32_INSTR_PT(328) OR ROM32_INSTR_PT(329)
     OR ROM32_INSTR_PT(332) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(337) OR ROM32_INSTR_PT(338)
     OR ROM32_INSTR_PT(339) OR ROM32_INSTR_PT(344)
     OR ROM32_INSTR_PT(346) OR ROM32_INSTR_PT(348)
     OR ROM32_INSTR_PT(350) OR ROM32_INSTR_PT(357)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(362)
     OR ROM32_INSTR_PT(363) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(368)
     OR ROM32_INSTR_PT(371) OR ROM32_INSTR_PT(373)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(378) OR ROM32_INSTR_PT(379)
     OR ROM32_INSTR_PT(381) OR ROM32_INSTR_PT(382)
     OR ROM32_INSTR_PT(383) OR ROM32_INSTR_PT(386)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(388)
     OR ROM32_INSTR_PT(390) OR ROM32_INSTR_PT(392)
     OR ROM32_INSTR_PT(393) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(395) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(400)
     OR ROM32_INSTR_PT(401) OR ROM32_INSTR_PT(402)
     OR ROM32_INSTR_PT(404) OR ROM32_INSTR_PT(405)
     OR ROM32_INSTR_PT(406) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(411) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(416)
     OR ROM32_INSTR_PT(417) OR ROM32_INSTR_PT(418)
     OR ROM32_INSTR_PT(419) OR ROM32_INSTR_PT(421)
     OR ROM32_INSTR_PT(422) OR ROM32_INSTR_PT(423)
     OR ROM32_INSTR_PT(424) OR ROM32_INSTR_PT(425)
     OR ROM32_INSTR_PT(426) OR ROM32_INSTR_PT(433)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(435)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(437)
     OR ROM32_INSTR_PT(438) OR ROM32_INSTR_PT(441)
     OR ROM32_INSTR_PT(442) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(446) OR ROM32_INSTR_PT(451)
     OR ROM32_INSTR_PT(452) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(456)
     OR ROM32_INSTR_PT(458) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(463) OR ROM32_INSTR_PT(464)
     OR ROM32_INSTR_PT(465) OR ROM32_INSTR_PT(467)
     OR ROM32_INSTR_PT(468) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(471) OR ROM32_INSTR_PT(472)
     OR ROM32_INSTR_PT(474) OR ROM32_INSTR_PT(475)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(480)
     OR ROM32_INSTR_PT(481) OR ROM32_INSTR_PT(482)
     OR ROM32_INSTR_PT(484) OR ROM32_INSTR_PT(486)
     OR ROM32_INSTR_PT(489) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(494) OR ROM32_INSTR_PT(495)
     OR ROM32_INSTR_PT(496) OR ROM32_INSTR_PT(497)
     OR ROM32_INSTR_PT(502) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(505) OR ROM32_INSTR_PT(506)
     OR ROM32_INSTR_PT(507) OR ROM32_INSTR_PT(508)
     OR ROM32_INSTR_PT(513) OR ROM32_INSTR_PT(514)
     OR ROM32_INSTR_PT(517) OR ROM32_INSTR_PT(519)
     OR ROM32_INSTR_PT(520) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(524)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(537) OR ROM32_INSTR_PT(539)
     OR ROM32_INSTR_PT(541) OR ROM32_INSTR_PT(544)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(549)
     OR ROM32_INSTR_PT(550) OR ROM32_INSTR_PT(551)
     OR ROM32_INSTR_PT(552) OR ROM32_INSTR_PT(554)
     OR ROM32_INSTR_PT(556) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(561)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(568)
     OR ROM32_INSTR_PT(569) OR ROM32_INSTR_PT(570)
     OR ROM32_INSTR_PT(571) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(575) OR ROM32_INSTR_PT(577)
     OR ROM32_INSTR_PT(578) OR ROM32_INSTR_PT(579)
     OR ROM32_INSTR_PT(580) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(582) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(584) OR ROM32_INSTR_PT(585)
     OR ROM32_INSTR_PT(586) OR ROM32_INSTR_PT(587)
     OR ROM32_INSTR_PT(588) OR ROM32_INSTR_PT(590)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(593)
     OR ROM32_INSTR_PT(595) OR ROM32_INSTR_PT(596)
     OR ROM32_INSTR_PT(598) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(602)
     OR ROM32_INSTR_PT(604) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(606) OR ROM32_INSTR_PT(607)
     OR ROM32_INSTR_PT(608) OR ROM32_INSTR_PT(609)
     OR ROM32_INSTR_PT(610) OR ROM32_INSTR_PT(611)
     OR ROM32_INSTR_PT(612) OR ROM32_INSTR_PT(614)
     OR ROM32_INSTR_PT(620) OR ROM32_INSTR_PT(621)
     OR ROM32_INSTR_PT(624) OR ROM32_INSTR_PT(625)
     OR ROM32_INSTR_PT(626) OR ROM32_INSTR_PT(629)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(632)
     OR ROM32_INSTR_PT(634) OR ROM32_INSTR_PT(638)
     OR ROM32_INSTR_PT(639) OR ROM32_INSTR_PT(640)
     OR ROM32_INSTR_PT(642) OR ROM32_INSTR_PT(643)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(653)
     OR ROM32_INSTR_PT(657) OR ROM32_INSTR_PT(659)
     OR ROM32_INSTR_PT(660) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(664) OR ROM32_INSTR_PT(666)
     OR ROM32_INSTR_PT(668) OR ROM32_INSTR_PT(672)
     OR ROM32_INSTR_PT(677) OR ROM32_INSTR_PT(680)
     OR ROM32_INSTR_PT(684) OR ROM32_INSTR_PT(689)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(698)
     OR ROM32_INSTR_PT(702) OR ROM32_INSTR_PT(704)
     OR ROM32_INSTR_PT(708) OR ROM32_INSTR_PT(713)
     OR ROM32_INSTR_PT(718) OR ROM32_INSTR_PT(719)
     OR ROM32_INSTR_PT(720) OR ROM32_INSTR_PT(726)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(729)
     OR ROM32_INSTR_PT(736) OR ROM32_INSTR_PT(751)
     OR ROM32_INSTR_PT(752) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(755) OR ROM32_INSTR_PT(759)
     OR ROM32_INSTR_PT(762) OR ROM32_INSTR_PT(770)
     OR ROM32_INSTR_PT(774) OR ROM32_INSTR_PT(787)
     OR ROM32_INSTR_PT(790) OR ROM32_INSTR_PT(792)
     OR ROM32_INSTR_PT(803) OR ROM32_INSTR_PT(805)
     OR ROM32_INSTR_PT(807) OR ROM32_INSTR_PT(812)
     OR ROM32_INSTR_PT(817) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(823) OR ROM32_INSTR_PT(831)
     OR ROM32_INSTR_PT(845) OR ROM32_INSTR_PT(853)
     OR ROM32_INSTR_PT(854) OR ROM32_INSTR_PT(855)
     OR ROM32_INSTR_PT(857) OR ROM32_INSTR_PT(862)
     OR ROM32_INSTR_PT(869) OR ROM32_INSTR_PT(870)
     OR ROM32_INSTR_PT(878) OR ROM32_INSTR_PT(881)
    );
MQQ1859:TEMPLATE(4) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(7)
     OR ROM32_INSTR_PT(13) OR ROM32_INSTR_PT(14)
     OR ROM32_INSTR_PT(18) OR ROM32_INSTR_PT(23)
     OR ROM32_INSTR_PT(27) OR ROM32_INSTR_PT(28)
     OR ROM32_INSTR_PT(29) OR ROM32_INSTR_PT(31)
     OR ROM32_INSTR_PT(33) OR ROM32_INSTR_PT(35)
     OR ROM32_INSTR_PT(38) OR ROM32_INSTR_PT(39)
     OR ROM32_INSTR_PT(41) OR ROM32_INSTR_PT(42)
     OR ROM32_INSTR_PT(43) OR ROM32_INSTR_PT(45)
     OR ROM32_INSTR_PT(53) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(62)
     OR ROM32_INSTR_PT(68) OR ROM32_INSTR_PT(70)
     OR ROM32_INSTR_PT(72) OR ROM32_INSTR_PT(76)
     OR ROM32_INSTR_PT(79) OR ROM32_INSTR_PT(80)
     OR ROM32_INSTR_PT(81) OR ROM32_INSTR_PT(83)
     OR ROM32_INSTR_PT(85) OR ROM32_INSTR_PT(92)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(98) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(102) OR ROM32_INSTR_PT(105)
     OR ROM32_INSTR_PT(109) OR ROM32_INSTR_PT(110)
     OR ROM32_INSTR_PT(111) OR ROM32_INSTR_PT(113)
     OR ROM32_INSTR_PT(117) OR ROM32_INSTR_PT(120)
     OR ROM32_INSTR_PT(122) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(128) OR ROM32_INSTR_PT(130)
     OR ROM32_INSTR_PT(138) OR ROM32_INSTR_PT(139)
     OR ROM32_INSTR_PT(141) OR ROM32_INSTR_PT(142)
     OR ROM32_INSTR_PT(144) OR ROM32_INSTR_PT(145)
     OR ROM32_INSTR_PT(146) OR ROM32_INSTR_PT(147)
     OR ROM32_INSTR_PT(150) OR ROM32_INSTR_PT(151)
     OR ROM32_INSTR_PT(153) OR ROM32_INSTR_PT(155)
     OR ROM32_INSTR_PT(158) OR ROM32_INSTR_PT(159)
     OR ROM32_INSTR_PT(162) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(165) OR ROM32_INSTR_PT(166)
     OR ROM32_INSTR_PT(172) OR ROM32_INSTR_PT(173)
     OR ROM32_INSTR_PT(174) OR ROM32_INSTR_PT(175)
     OR ROM32_INSTR_PT(176) OR ROM32_INSTR_PT(177)
     OR ROM32_INSTR_PT(178) OR ROM32_INSTR_PT(180)
     OR ROM32_INSTR_PT(181) OR ROM32_INSTR_PT(185)
     OR ROM32_INSTR_PT(186) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(189) OR ROM32_INSTR_PT(192)
     OR ROM32_INSTR_PT(193) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(199) OR ROM32_INSTR_PT(203)
     OR ROM32_INSTR_PT(205) OR ROM32_INSTR_PT(206)
     OR ROM32_INSTR_PT(207) OR ROM32_INSTR_PT(208)
     OR ROM32_INSTR_PT(209) OR ROM32_INSTR_PT(210)
     OR ROM32_INSTR_PT(212) OR ROM32_INSTR_PT(218)
     OR ROM32_INSTR_PT(222) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(228) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(230) OR ROM32_INSTR_PT(232)
     OR ROM32_INSTR_PT(233) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(237) OR ROM32_INSTR_PT(240)
     OR ROM32_INSTR_PT(242) OR ROM32_INSTR_PT(245)
     OR ROM32_INSTR_PT(249) OR ROM32_INSTR_PT(251)
     OR ROM32_INSTR_PT(252) OR ROM32_INSTR_PT(254)
     OR ROM32_INSTR_PT(255) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(262)
     OR ROM32_INSTR_PT(266) OR ROM32_INSTR_PT(268)
     OR ROM32_INSTR_PT(272) OR ROM32_INSTR_PT(275)
     OR ROM32_INSTR_PT(279) OR ROM32_INSTR_PT(285)
     OR ROM32_INSTR_PT(287) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(290) OR ROM32_INSTR_PT(291)
     OR ROM32_INSTR_PT(292) OR ROM32_INSTR_PT(294)
     OR ROM32_INSTR_PT(302) OR ROM32_INSTR_PT(305)
     OR ROM32_INSTR_PT(307) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(311) OR ROM32_INSTR_PT(318)
     OR ROM32_INSTR_PT(322) OR ROM32_INSTR_PT(323)
     OR ROM32_INSTR_PT(325) OR ROM32_INSTR_PT(329)
     OR ROM32_INSTR_PT(332) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(337) OR ROM32_INSTR_PT(338)
     OR ROM32_INSTR_PT(339) OR ROM32_INSTR_PT(344)
     OR ROM32_INSTR_PT(346) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(356) OR ROM32_INSTR_PT(357)
     OR ROM32_INSTR_PT(358) OR ROM32_INSTR_PT(359)
     OR ROM32_INSTR_PT(362) OR ROM32_INSTR_PT(363)
     OR ROM32_INSTR_PT(365) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(368)
     OR ROM32_INSTR_PT(370) OR ROM32_INSTR_PT(373)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(378) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(382) OR ROM32_INSTR_PT(386)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(388)
     OR ROM32_INSTR_PT(391) OR ROM32_INSTR_PT(393)
     OR ROM32_INSTR_PT(394) OR ROM32_INSTR_PT(395)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(399)
     OR ROM32_INSTR_PT(400) OR ROM32_INSTR_PT(402)
     OR ROM32_INSTR_PT(404) OR ROM32_INSTR_PT(405)
     OR ROM32_INSTR_PT(409) OR ROM32_INSTR_PT(415)
     OR ROM32_INSTR_PT(416) OR ROM32_INSTR_PT(417)
     OR ROM32_INSTR_PT(418) OR ROM32_INSTR_PT(419)
     OR ROM32_INSTR_PT(422) OR ROM32_INSTR_PT(423)
     OR ROM32_INSTR_PT(425) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(435)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(438)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(442)
     OR ROM32_INSTR_PT(443) OR ROM32_INSTR_PT(446)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(452)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(456)
     OR ROM32_INSTR_PT(458) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(463) OR ROM32_INSTR_PT(464)
     OR ROM32_INSTR_PT(465) OR ROM32_INSTR_PT(467)
     OR ROM32_INSTR_PT(468) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(471) OR ROM32_INSTR_PT(472)
     OR ROM32_INSTR_PT(473) OR ROM32_INSTR_PT(474)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(480)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(489)
     OR ROM32_INSTR_PT(496) OR ROM32_INSTR_PT(497)
     OR ROM32_INSTR_PT(498) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(505) OR ROM32_INSTR_PT(507)
     OR ROM32_INSTR_PT(513) OR ROM32_INSTR_PT(514)
     OR ROM32_INSTR_PT(517) OR ROM32_INSTR_PT(527)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(537)
     OR ROM32_INSTR_PT(539) OR ROM32_INSTR_PT(541)
     OR ROM32_INSTR_PT(544) OR ROM32_INSTR_PT(547)
     OR ROM32_INSTR_PT(549) OR ROM32_INSTR_PT(551)
     OR ROM32_INSTR_PT(555) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(561)
     OR ROM32_INSTR_PT(563) OR ROM32_INSTR_PT(566)
     OR ROM32_INSTR_PT(569) OR ROM32_INSTR_PT(570)
     OR ROM32_INSTR_PT(571) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(577) OR ROM32_INSTR_PT(579)
     OR ROM32_INSTR_PT(580) OR ROM32_INSTR_PT(584)
     OR ROM32_INSTR_PT(586) OR ROM32_INSTR_PT(587)
     OR ROM32_INSTR_PT(589) OR ROM32_INSTR_PT(591)
     OR ROM32_INSTR_PT(593) OR ROM32_INSTR_PT(596)
     OR ROM32_INSTR_PT(597) OR ROM32_INSTR_PT(598)
     OR ROM32_INSTR_PT(599) OR ROM32_INSTR_PT(600)
     OR ROM32_INSTR_PT(604) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(606) OR ROM32_INSTR_PT(607)
     OR ROM32_INSTR_PT(608) OR ROM32_INSTR_PT(609)
     OR ROM32_INSTR_PT(610) OR ROM32_INSTR_PT(611)
     OR ROM32_INSTR_PT(614) OR ROM32_INSTR_PT(620)
     OR ROM32_INSTR_PT(624) OR ROM32_INSTR_PT(625)
     OR ROM32_INSTR_PT(629) OR ROM32_INSTR_PT(632)
     OR ROM32_INSTR_PT(634) OR ROM32_INSTR_PT(638)
     OR ROM32_INSTR_PT(640) OR ROM32_INSTR_PT(641)
     OR ROM32_INSTR_PT(643) OR ROM32_INSTR_PT(652)
     OR ROM32_INSTR_PT(653) OR ROM32_INSTR_PT(659)
     OR ROM32_INSTR_PT(660) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(664) OR ROM32_INSTR_PT(668)
     OR ROM32_INSTR_PT(672) OR ROM32_INSTR_PT(680)
     OR ROM32_INSTR_PT(683) OR ROM32_INSTR_PT(684)
     OR ROM32_INSTR_PT(689) OR ROM32_INSTR_PT(691)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(697)
     OR ROM32_INSTR_PT(698) OR ROM32_INSTR_PT(702)
     OR ROM32_INSTR_PT(704) OR ROM32_INSTR_PT(708)
     OR ROM32_INSTR_PT(711) OR ROM32_INSTR_PT(713)
     OR ROM32_INSTR_PT(718) OR ROM32_INSTR_PT(720)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(729)
     OR ROM32_INSTR_PT(733) OR ROM32_INSTR_PT(751)
     OR ROM32_INSTR_PT(752) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(759) OR ROM32_INSTR_PT(763)
     OR ROM32_INSTR_PT(774) OR ROM32_INSTR_PT(787)
     OR ROM32_INSTR_PT(790) OR ROM32_INSTR_PT(792)
     OR ROM32_INSTR_PT(795) OR ROM32_INSTR_PT(801)
     OR ROM32_INSTR_PT(803) OR ROM32_INSTR_PT(805)
     OR ROM32_INSTR_PT(807) OR ROM32_INSTR_PT(812)
     OR ROM32_INSTR_PT(817) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(823) OR ROM32_INSTR_PT(829)
     OR ROM32_INSTR_PT(831) OR ROM32_INSTR_PT(845)
     OR ROM32_INSTR_PT(847) OR ROM32_INSTR_PT(851)
     OR ROM32_INSTR_PT(853) OR ROM32_INSTR_PT(854)
     OR ROM32_INSTR_PT(857) OR ROM32_INSTR_PT(869)
     OR ROM32_INSTR_PT(872) OR ROM32_INSTR_PT(878)
     OR ROM32_INSTR_PT(881));
MQQ1860:TEMPLATE(5) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(7)
     OR ROM32_INSTR_PT(9) OR ROM32_INSTR_PT(10)
     OR ROM32_INSTR_PT(12) OR ROM32_INSTR_PT(13)
     OR ROM32_INSTR_PT(14) OR ROM32_INSTR_PT(20)
     OR ROM32_INSTR_PT(26) OR ROM32_INSTR_PT(33)
     OR ROM32_INSTR_PT(37) OR ROM32_INSTR_PT(39)
     OR ROM32_INSTR_PT(41) OR ROM32_INSTR_PT(42)
     OR ROM32_INSTR_PT(45) OR ROM32_INSTR_PT(49)
     OR ROM32_INSTR_PT(51) OR ROM32_INSTR_PT(52)
     OR ROM32_INSTR_PT(53) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(59)
     OR ROM32_INSTR_PT(63) OR ROM32_INSTR_PT(66)
     OR ROM32_INSTR_PT(67) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(73) OR ROM32_INSTR_PT(83)
     OR ROM32_INSTR_PT(84) OR ROM32_INSTR_PT(85)
     OR ROM32_INSTR_PT(87) OR ROM32_INSTR_PT(90)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(96)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(102) OR ROM32_INSTR_PT(103)
     OR ROM32_INSTR_PT(106) OR ROM32_INSTR_PT(109)
     OR ROM32_INSTR_PT(110) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(124) OR ROM32_INSTR_PT(130)
     OR ROM32_INSTR_PT(131) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(139) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(142) OR ROM32_INSTR_PT(143)
     OR ROM32_INSTR_PT(144) OR ROM32_INSTR_PT(153)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(159) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(164) OR ROM32_INSTR_PT(169)
     OR ROM32_INSTR_PT(170) OR ROM32_INSTR_PT(176)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(180)
     OR ROM32_INSTR_PT(181) OR ROM32_INSTR_PT(183)
     OR ROM32_INSTR_PT(184) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(192) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(196) OR ROM32_INSTR_PT(199)
     OR ROM32_INSTR_PT(202) OR ROM32_INSTR_PT(203)
     OR ROM32_INSTR_PT(204) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(206) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(212) OR ROM32_INSTR_PT(216)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(232)
     OR ROM32_INSTR_PT(233) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(241)
     OR ROM32_INSTR_PT(243) OR ROM32_INSTR_PT(244)
     OR ROM32_INSTR_PT(249) OR ROM32_INSTR_PT(252)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(259) OR ROM32_INSTR_PT(260)
     OR ROM32_INSTR_PT(261) OR ROM32_INSTR_PT(264)
     OR ROM32_INSTR_PT(266) OR ROM32_INSTR_PT(267)
     OR ROM32_INSTR_PT(268) OR ROM32_INSTR_PT(269)
     OR ROM32_INSTR_PT(271) OR ROM32_INSTR_PT(274)
     OR ROM32_INSTR_PT(276) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(280) OR ROM32_INSTR_PT(282)
     OR ROM32_INSTR_PT(284) OR ROM32_INSTR_PT(288)
     OR ROM32_INSTR_PT(290) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(306) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(310) OR ROM32_INSTR_PT(318)
     OR ROM32_INSTR_PT(323) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(346)
     OR ROM32_INSTR_PT(348) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(353) OR ROM32_INSTR_PT(356)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(363)
     OR ROM32_INSTR_PT(364) OR ROM32_INSTR_PT(367)
     OR ROM32_INSTR_PT(371) OR ROM32_INSTR_PT(373)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(382) OR ROM32_INSTR_PT(383)
     OR ROM32_INSTR_PT(386) OR ROM32_INSTR_PT(390)
     OR ROM32_INSTR_PT(392) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(396) OR ROM32_INSTR_PT(400)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(405)
     OR ROM32_INSTR_PT(406) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(413) OR ROM32_INSTR_PT(415)
     OR ROM32_INSTR_PT(417) OR ROM32_INSTR_PT(422)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(425) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(428) OR ROM32_INSTR_PT(430)
     OR ROM32_INSTR_PT(431) OR ROM32_INSTR_PT(434)
     OR ROM32_INSTR_PT(435) OR ROM32_INSTR_PT(436)
     OR ROM32_INSTR_PT(438) OR ROM32_INSTR_PT(441)
     OR ROM32_INSTR_PT(442) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(445) OR ROM32_INSTR_PT(449)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(452)
     OR ROM32_INSTR_PT(453) OR ROM32_INSTR_PT(458)
     OR ROM32_INSTR_PT(464) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(474)
     OR ROM32_INSTR_PT(475) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(481)
     OR ROM32_INSTR_PT(482) OR ROM32_INSTR_PT(484)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(491) OR ROM32_INSTR_PT(494)
     OR ROM32_INSTR_PT(495) OR ROM32_INSTR_PT(501)
     OR ROM32_INSTR_PT(503) OR ROM32_INSTR_PT(507)
     OR ROM32_INSTR_PT(509) OR ROM32_INSTR_PT(511)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(517)
     OR ROM32_INSTR_PT(520) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(524)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(531)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(541) OR ROM32_INSTR_PT(544)
     OR ROM32_INSTR_PT(550) OR ROM32_INSTR_PT(551)
     OR ROM32_INSTR_PT(552) OR ROM32_INSTR_PT(554)
     OR ROM32_INSTR_PT(555) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(569)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(575)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(580)
     OR ROM32_INSTR_PT(581) OR ROM32_INSTR_PT(582)
     OR ROM32_INSTR_PT(583) OR ROM32_INSTR_PT(584)
     OR ROM32_INSTR_PT(588) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(601)
     OR ROM32_INSTR_PT(602) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(609) OR ROM32_INSTR_PT(610)
     OR ROM32_INSTR_PT(613) OR ROM32_INSTR_PT(615)
     OR ROM32_INSTR_PT(616) OR ROM32_INSTR_PT(617)
     OR ROM32_INSTR_PT(620) OR ROM32_INSTR_PT(622)
     OR ROM32_INSTR_PT(624) OR ROM32_INSTR_PT(626)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(634)
     OR ROM32_INSTR_PT(638) OR ROM32_INSTR_PT(639)
     OR ROM32_INSTR_PT(642) OR ROM32_INSTR_PT(643)
     OR ROM32_INSTR_PT(654) OR ROM32_INSTR_PT(660)
     OR ROM32_INSTR_PT(663) OR ROM32_INSTR_PT(664)
     OR ROM32_INSTR_PT(666) OR ROM32_INSTR_PT(674)
     OR ROM32_INSTR_PT(677) OR ROM32_INSTR_PT(684)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(693)
     OR ROM32_INSTR_PT(697) OR ROM32_INSTR_PT(708)
     OR ROM32_INSTR_PT(711) OR ROM32_INSTR_PT(713)
     OR ROM32_INSTR_PT(718) OR ROM32_INSTR_PT(719)
     OR ROM32_INSTR_PT(726) OR ROM32_INSTR_PT(729)
     OR ROM32_INSTR_PT(745) OR ROM32_INSTR_PT(755)
     OR ROM32_INSTR_PT(762) OR ROM32_INSTR_PT(763)
     OR ROM32_INSTR_PT(792) OR ROM32_INSTR_PT(805)
     OR ROM32_INSTR_PT(812) OR ROM32_INSTR_PT(818)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(829)
     OR ROM32_INSTR_PT(831) OR ROM32_INSTR_PT(845)
     OR ROM32_INSTR_PT(853) OR ROM32_INSTR_PT(854)
     OR ROM32_INSTR_PT(855) OR ROM32_INSTR_PT(857)
     OR ROM32_INSTR_PT(862) OR ROM32_INSTR_PT(870)
     OR ROM32_INSTR_PT(872) OR ROM32_INSTR_PT(878)
    );
MQQ1861:TEMPLATE(6) <= 
    ('0');
MQQ1862:TEMPLATE(7) <= 
    ('0');
MQQ1863:TEMPLATE(8) <= 
    ('0');
MQQ1864:TEMPLATE(9) <= 
    (ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(8)
     OR ROM32_INSTR_PT(10) OR ROM32_INSTR_PT(12)
     OR ROM32_INSTR_PT(14) OR ROM32_INSTR_PT(17)
     OR ROM32_INSTR_PT(23) OR ROM32_INSTR_PT(28)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(37)
     OR ROM32_INSTR_PT(42) OR ROM32_INSTR_PT(45)
     OR ROM32_INSTR_PT(53) OR ROM32_INSTR_PT(55)
     OR ROM32_INSTR_PT(56) OR ROM32_INSTR_PT(60)
     OR ROM32_INSTR_PT(63) OR ROM32_INSTR_PT(73)
     OR ROM32_INSTR_PT(74) OR ROM32_INSTR_PT(85)
     OR ROM32_INSTR_PT(87) OR ROM32_INSTR_PT(90)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(102)
     OR ROM32_INSTR_PT(103) OR ROM32_INSTR_PT(105)
     OR ROM32_INSTR_PT(106) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(120) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(130) OR ROM32_INSTR_PT(134)
     OR ROM32_INSTR_PT(135) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(142) OR ROM32_INSTR_PT(148)
     OR ROM32_INSTR_PT(154) OR ROM32_INSTR_PT(155)
     OR ROM32_INSTR_PT(162) OR ROM32_INSTR_PT(172)
     OR ROM32_INSTR_PT(174) OR ROM32_INSTR_PT(175)
     OR ROM32_INSTR_PT(176) OR ROM32_INSTR_PT(177)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(180)
     OR ROM32_INSTR_PT(181) OR ROM32_INSTR_PT(184)
     OR ROM32_INSTR_PT(187) OR ROM32_INSTR_PT(192)
     OR ROM32_INSTR_PT(193) OR ROM32_INSTR_PT(199)
     OR ROM32_INSTR_PT(202) OR ROM32_INSTR_PT(209)
     OR ROM32_INSTR_PT(214) OR ROM32_INSTR_PT(216)
     OR ROM32_INSTR_PT(218) OR ROM32_INSTR_PT(222)
     OR ROM32_INSTR_PT(223) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(232)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(240)
     OR ROM32_INSTR_PT(242) OR ROM32_INSTR_PT(244)
     OR ROM32_INSTR_PT(249) OR ROM32_INSTR_PT(255)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(258)
     OR ROM32_INSTR_PT(260) OR ROM32_INSTR_PT(269)
     OR ROM32_INSTR_PT(272) OR ROM32_INSTR_PT(273)
     OR ROM32_INSTR_PT(274) OR ROM32_INSTR_PT(275)
     OR ROM32_INSTR_PT(280) OR ROM32_INSTR_PT(282)
     OR ROM32_INSTR_PT(283) OR ROM32_INSTR_PT(287)
     OR ROM32_INSTR_PT(288) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(297)
     OR ROM32_INSTR_PT(299) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(309) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(319)
     OR ROM32_INSTR_PT(321) OR ROM32_INSTR_PT(338)
     OR ROM32_INSTR_PT(345) OR ROM32_INSTR_PT(348)
     OR ROM32_INSTR_PT(353) OR ROM32_INSTR_PT(357)
     OR ROM32_INSTR_PT(359) OR ROM32_INSTR_PT(362)
     OR ROM32_INSTR_PT(363) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(374)
     OR ROM32_INSTR_PT(377) OR ROM32_INSTR_PT(378)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(382)
     OR ROM32_INSTR_PT(383) OR ROM32_INSTR_PT(386)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(388)
     OR ROM32_INSTR_PT(391) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(395) OR ROM32_INSTR_PT(399)
     OR ROM32_INSTR_PT(400) OR ROM32_INSTR_PT(401)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(406)
     OR ROM32_INSTR_PT(409) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(416)
     OR ROM32_INSTR_PT(422) OR ROM32_INSTR_PT(423)
     OR ROM32_INSTR_PT(431) OR ROM32_INSTR_PT(433)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(436)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(464) OR ROM32_INSTR_PT(467)
     OR ROM32_INSTR_PT(469) OR ROM32_INSTR_PT(471)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(475)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(482)
     OR ROM32_INSTR_PT(489) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(491) OR ROM32_INSTR_PT(494)
     OR ROM32_INSTR_PT(497) OR ROM32_INSTR_PT(498)
     OR ROM32_INSTR_PT(501) OR ROM32_INSTR_PT(502)
     OR ROM32_INSTR_PT(504) OR ROM32_INSTR_PT(506)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(516)
     OR ROM32_INSTR_PT(517) OR ROM32_INSTR_PT(519)
     OR ROM32_INSTR_PT(520) OR ROM32_INSTR_PT(532)
     OR ROM32_INSTR_PT(534) OR ROM32_INSTR_PT(535)
     OR ROM32_INSTR_PT(543) OR ROM32_INSTR_PT(544)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(550)
     OR ROM32_INSTR_PT(552) OR ROM32_INSTR_PT(556)
     OR ROM32_INSTR_PT(557) OR ROM32_INSTR_PT(568)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(571)
     OR ROM32_INSTR_PT(574) OR ROM32_INSTR_PT(575)
     OR ROM32_INSTR_PT(586) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(589) OR ROM32_INSTR_PT(590)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(602)
     OR ROM32_INSTR_PT(604) OR ROM32_INSTR_PT(606)
     OR ROM32_INSTR_PT(609) OR ROM32_INSTR_PT(611)
     OR ROM32_INSTR_PT(612) OR ROM32_INSTR_PT(613)
     OR ROM32_INSTR_PT(621) OR ROM32_INSTR_PT(625)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(639)
     OR ROM32_INSTR_PT(640) OR ROM32_INSTR_PT(646)
     OR ROM32_INSTR_PT(647) OR ROM32_INSTR_PT(652)
     OR ROM32_INSTR_PT(659) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(666) OR ROM32_INSTR_PT(677)
     OR ROM32_INSTR_PT(689) OR ROM32_INSTR_PT(690)
     OR ROM32_INSTR_PT(698) OR ROM32_INSTR_PT(700)
     OR ROM32_INSTR_PT(733) OR ROM32_INSTR_PT(745)
     OR ROM32_INSTR_PT(751) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(790) OR ROM32_INSTR_PT(807)
     OR ROM32_INSTR_PT(823) OR ROM32_INSTR_PT(845)
    );
MQQ1865:TEMPLATE(10) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(13)
     OR ROM32_INSTR_PT(14) OR ROM32_INSTR_PT(16)
     OR ROM32_INSTR_PT(18) OR ROM32_INSTR_PT(32)
     OR ROM32_INSTR_PT(38) OR ROM32_INSTR_PT(41)
     OR ROM32_INSTR_PT(42) OR ROM32_INSTR_PT(45)
     OR ROM32_INSTR_PT(51) OR ROM32_INSTR_PT(52)
     OR ROM32_INSTR_PT(53) OR ROM32_INSTR_PT(57)
     OR ROM32_INSTR_PT(76) OR ROM32_INSTR_PT(77)
     OR ROM32_INSTR_PT(85) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(99) OR ROM32_INSTR_PT(113)
     OR ROM32_INSTR_PT(114) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(123)
     OR ROM32_INSTR_PT(125) OR ROM32_INSTR_PT(127)
     OR ROM32_INSTR_PT(128) OR ROM32_INSTR_PT(130)
     OR ROM32_INSTR_PT(138) OR ROM32_INSTR_PT(139)
     OR ROM32_INSTR_PT(142) OR ROM32_INSTR_PT(143)
     OR ROM32_INSTR_PT(153) OR ROM32_INSTR_PT(169)
     OR ROM32_INSTR_PT(171) OR ROM32_INSTR_PT(173)
     OR ROM32_INSTR_PT(174) OR ROM32_INSTR_PT(180)
     OR ROM32_INSTR_PT(181) OR ROM32_INSTR_PT(183)
     OR ROM32_INSTR_PT(189) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(200) OR ROM32_INSTR_PT(203)
     OR ROM32_INSTR_PT(204) OR ROM32_INSTR_PT(214)
     OR ROM32_INSTR_PT(219) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(235) OR ROM32_INSTR_PT(237)
     OR ROM32_INSTR_PT(240) OR ROM32_INSTR_PT(241)
     OR ROM32_INSTR_PT(250) OR ROM32_INSTR_PT(251)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(261) OR ROM32_INSTR_PT(267)
     OR ROM32_INSTR_PT(270) OR ROM32_INSTR_PT(271)
     OR ROM32_INSTR_PT(274) OR ROM32_INSTR_PT(276)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(328) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(363)
     OR ROM32_INSTR_PT(364) OR ROM32_INSTR_PT(365)
     OR ROM32_INSTR_PT(370) OR ROM32_INSTR_PT(371)
     OR ROM32_INSTR_PT(376) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(390) OR ROM32_INSTR_PT(395)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(400)
     OR ROM32_INSTR_PT(404) OR ROM32_INSTR_PT(418)
     OR ROM32_INSTR_PT(419) OR ROM32_INSTR_PT(421)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(439)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(446)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(468)
     OR ROM32_INSTR_PT(473) OR ROM32_INSTR_PT(477)
     OR ROM32_INSTR_PT(478) OR ROM32_INSTR_PT(480)
     OR ROM32_INSTR_PT(489) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(504) OR ROM32_INSTR_PT(505)
     OR ROM32_INSTR_PT(508) OR ROM32_INSTR_PT(509)
     OR ROM32_INSTR_PT(517) OR ROM32_INSTR_PT(524)
     OR ROM32_INSTR_PT(527) OR ROM32_INSTR_PT(531)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(537)
     OR ROM32_INSTR_PT(538) OR ROM32_INSTR_PT(546)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(555)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(562)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(578)
     OR ROM32_INSTR_PT(582) OR ROM32_INSTR_PT(585)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(593)
     OR ROM32_INSTR_PT(595) OR ROM32_INSTR_PT(597)
     OR ROM32_INSTR_PT(598) OR ROM32_INSTR_PT(603)
     OR ROM32_INSTR_PT(608) OR ROM32_INSTR_PT(615)
     OR ROM32_INSTR_PT(624) OR ROM32_INSTR_PT(626)
     OR ROM32_INSTR_PT(629) OR ROM32_INSTR_PT(635)
     OR ROM32_INSTR_PT(641) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(654)
     OR ROM32_INSTR_PT(680) OR ROM32_INSTR_PT(683)
     OR ROM32_INSTR_PT(689) OR ROM32_INSTR_PT(708)
     OR ROM32_INSTR_PT(713) OR ROM32_INSTR_PT(718)
     OR ROM32_INSTR_PT(720) OR ROM32_INSTR_PT(728)
     OR ROM32_INSTR_PT(729) OR ROM32_INSTR_PT(731)
     OR ROM32_INSTR_PT(755) OR ROM32_INSTR_PT(763)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(857)
     OR ROM32_INSTR_PT(872));
MQQ1866:TEMPLATE(11) <= 
    ('0');
MQQ1867:TEMPLATE(12) <= 
    ('0');
MQQ1868:TEMPLATE(13) <= 
    ('0');
MQQ1869:TEMPLATE(14) <= 
    (ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(10)
     OR ROM32_INSTR_PT(12) OR ROM32_INSTR_PT(14)
     OR ROM32_INSTR_PT(16) OR ROM32_INSTR_PT(20)
     OR ROM32_INSTR_PT(23) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(32) OR ROM32_INSTR_PT(34)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(37)
     OR ROM32_INSTR_PT(42) OR ROM32_INSTR_PT(52)
     OR ROM32_INSTR_PT(53) OR ROM32_INSTR_PT(55)
     OR ROM32_INSTR_PT(56) OR ROM32_INSTR_PT(63)
     OR ROM32_INSTR_PT(67) OR ROM32_INSTR_PT(73)
     OR ROM32_INSTR_PT(77) OR ROM32_INSTR_PT(79)
     OR ROM32_INSTR_PT(85) OR ROM32_INSTR_PT(87)
     OR ROM32_INSTR_PT(90) OR ROM32_INSTR_PT(92)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(99) OR ROM32_INSTR_PT(103)
     OR ROM32_INSTR_PT(105) OR ROM32_INSTR_PT(111)
     OR ROM32_INSTR_PT(114) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(125) OR ROM32_INSTR_PT(127)
     OR ROM32_INSTR_PT(130) OR ROM32_INSTR_PT(138)
     OR ROM32_INSTR_PT(143) OR ROM32_INSTR_PT(155)
     OR ROM32_INSTR_PT(169) OR ROM32_INSTR_PT(171)
     OR ROM32_INSTR_PT(172) OR ROM32_INSTR_PT(174)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(181)
     OR ROM32_INSTR_PT(184) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(196) OR ROM32_INSTR_PT(200)
     OR ROM32_INSTR_PT(202) OR ROM32_INSTR_PT(209)
     OR ROM32_INSTR_PT(214) OR ROM32_INSTR_PT(216)
     OR ROM32_INSTR_PT(218) OR ROM32_INSTR_PT(219)
     OR ROM32_INSTR_PT(224) OR ROM32_INSTR_PT(227)
     OR ROM32_INSTR_PT(229) OR ROM32_INSTR_PT(232)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(240)
     OR ROM32_INSTR_PT(250) OR ROM32_INSTR_PT(257)
     OR ROM32_INSTR_PT(259) OR ROM32_INSTR_PT(261)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(267)
     OR ROM32_INSTR_PT(269) OR ROM32_INSTR_PT(270)
     OR ROM32_INSTR_PT(271) OR ROM32_INSTR_PT(272)
     OR ROM32_INSTR_PT(273) OR ROM32_INSTR_PT(274)
     OR ROM32_INSTR_PT(275) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(280) OR ROM32_INSTR_PT(283)
     OR ROM32_INSTR_PT(284) OR ROM32_INSTR_PT(288)
     OR ROM32_INSTR_PT(290) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(299) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(309) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(321) OR ROM32_INSTR_PT(328)
     OR ROM32_INSTR_PT(345) OR ROM32_INSTR_PT(348)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(362)
     OR ROM32_INSTR_PT(363) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(368)
     OR ROM32_INSTR_PT(370) OR ROM32_INSTR_PT(371)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(383)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(390)
     OR ROM32_INSTR_PT(392) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(395) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(400) OR ROM32_INSTR_PT(401)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(406)
     OR ROM32_INSTR_PT(411) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(418) OR ROM32_INSTR_PT(421)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(433) OR ROM32_INSTR_PT(436)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(445)
     OR ROM32_INSTR_PT(449) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(456) OR ROM32_INSTR_PT(464)
     OR ROM32_INSTR_PT(469) OR ROM32_INSTR_PT(472)
     OR ROM32_INSTR_PT(475) OR ROM32_INSTR_PT(476)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(480)
     OR ROM32_INSTR_PT(481) OR ROM32_INSTR_PT(482)
     OR ROM32_INSTR_PT(484) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(494) OR ROM32_INSTR_PT(497)
     OR ROM32_INSTR_PT(502) OR ROM32_INSTR_PT(508)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(517)
     OR ROM32_INSTR_PT(519) OR ROM32_INSTR_PT(520)
     OR ROM32_INSTR_PT(521) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(524) OR ROM32_INSTR_PT(532)
     OR ROM32_INSTR_PT(534) OR ROM32_INSTR_PT(535)
     OR ROM32_INSTR_PT(536) OR ROM32_INSTR_PT(541)
     OR ROM32_INSTR_PT(543) OR ROM32_INSTR_PT(546)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(550)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(556)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(565)
     OR ROM32_INSTR_PT(568) OR ROM32_INSTR_PT(570)
     OR ROM32_INSTR_PT(574) OR ROM32_INSTR_PT(575)
     OR ROM32_INSTR_PT(578) OR ROM32_INSTR_PT(582)
     OR ROM32_INSTR_PT(585) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(590) OR ROM32_INSTR_PT(595)
     OR ROM32_INSTR_PT(602) OR ROM32_INSTR_PT(603)
     OR ROM32_INSTR_PT(606) OR ROM32_INSTR_PT(607)
     OR ROM32_INSTR_PT(611) OR ROM32_INSTR_PT(612)
     OR ROM32_INSTR_PT(617) OR ROM32_INSTR_PT(621)
     OR ROM32_INSTR_PT(625) OR ROM32_INSTR_PT(630)
     OR ROM32_INSTR_PT(633) OR ROM32_INSTR_PT(635)
     OR ROM32_INSTR_PT(639) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(647)
     OR ROM32_INSTR_PT(666) OR ROM32_INSTR_PT(677)
     OR ROM32_INSTR_PT(680) OR ROM32_INSTR_PT(689)
     OR ROM32_INSTR_PT(690) OR ROM32_INSTR_PT(698)
     OR ROM32_INSTR_PT(718) OR ROM32_INSTR_PT(731)
     OR ROM32_INSTR_PT(736) OR ROM32_INSTR_PT(745)
     OR ROM32_INSTR_PT(755) OR ROM32_INSTR_PT(762)
     OR ROM32_INSTR_PT(770) OR ROM32_INSTR_PT(818)
     OR ROM32_INSTR_PT(855) OR ROM32_INSTR_PT(862)
     OR ROM32_INSTR_PT(870));
MQQ1870:TEMPLATE(15) <= 
    (ROM32_INSTR_PT(8) OR ROM32_INSTR_PT(14)
     OR ROM32_INSTR_PT(17) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(34) OR ROM32_INSTR_PT(53)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(74)
     OR ROM32_INSTR_PT(79) OR ROM32_INSTR_PT(84)
     OR ROM32_INSTR_PT(92) OR ROM32_INSTR_PT(102)
     OR ROM32_INSTR_PT(111) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(117) OR ROM32_INSTR_PT(122)
     OR ROM32_INSTR_PT(123) OR ROM32_INSTR_PT(134)
     OR ROM32_INSTR_PT(141) OR ROM32_INSTR_PT(148)
     OR ROM32_INSTR_PT(159) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(170) OR ROM32_INSTR_PT(173)
     OR ROM32_INSTR_PT(174) OR ROM32_INSTR_PT(203)
     OR ROM32_INSTR_PT(212) OR ROM32_INSTR_PT(214)
     OR ROM32_INSTR_PT(215) OR ROM32_INSTR_PT(220)
     OR ROM32_INSTR_PT(223) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(240) OR ROM32_INSTR_PT(259)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(271)
     OR ROM32_INSTR_PT(276) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(290) OR ROM32_INSTR_PT(294)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(301)
     OR ROM32_INSTR_PT(309) OR ROM32_INSTR_PT(346)
     OR ROM32_INSTR_PT(350) OR ROM32_INSTR_PT(356)
     OR ROM32_INSTR_PT(360) OR ROM32_INSTR_PT(368)
     OR ROM32_INSTR_PT(376) OR ROM32_INSTR_PT(382)
     OR ROM32_INSTR_PT(386) OR ROM32_INSTR_PT(392)
     OR ROM32_INSTR_PT(395) OR ROM32_INSTR_PT(404)
     OR ROM32_INSTR_PT(413) OR ROM32_INSTR_PT(422)
     OR ROM32_INSTR_PT(430) OR ROM32_INSTR_PT(431)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(438)
     OR ROM32_INSTR_PT(439) OR ROM32_INSTR_PT(442)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(459)
     OR ROM32_INSTR_PT(471) OR ROM32_INSTR_PT(474)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(477)
     OR ROM32_INSTR_PT(503) OR ROM32_INSTR_PT(505)
     OR ROM32_INSTR_PT(506) OR ROM32_INSTR_PT(517)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(532)
     OR ROM32_INSTR_PT(536) OR ROM32_INSTR_PT(538)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(580) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(593) OR ROM32_INSTR_PT(598)
     OR ROM32_INSTR_PT(599) OR ROM32_INSTR_PT(607)
     OR ROM32_INSTR_PT(608) OR ROM32_INSTR_PT(620)
     OR ROM32_INSTR_PT(659) OR ROM32_INSTR_PT(664)
     OR ROM32_INSTR_PT(689) OR ROM32_INSTR_PT(692)
     OR ROM32_INSTR_PT(711) OR ROM32_INSTR_PT(726)
     OR ROM32_INSTR_PT(829) OR ROM32_INSTR_PT(831)
     OR ROM32_INSTR_PT(845) OR ROM32_INSTR_PT(853)
    );
MQQ1871:TEMPLATE(16) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(9)
     OR ROM32_INSTR_PT(16) OR ROM32_INSTR_PT(18)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(32) OR ROM32_INSTR_PT(34)
     OR ROM32_INSTR_PT(38) OR ROM32_INSTR_PT(49)
     OR ROM32_INSTR_PT(55) OR ROM32_INSTR_PT(67)
     OR ROM32_INSTR_PT(77) OR ROM32_INSTR_PT(79)
     OR ROM32_INSTR_PT(84) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(99) OR ROM32_INSTR_PT(105)
     OR ROM32_INSTR_PT(111) OR ROM32_INSTR_PT(114)
     OR ROM32_INSTR_PT(115) OR ROM32_INSTR_PT(118)
     OR ROM32_INSTR_PT(119) OR ROM32_INSTR_PT(122)
     OR ROM32_INSTR_PT(127) OR ROM32_INSTR_PT(171)
     OR ROM32_INSTR_PT(186) OR ROM32_INSTR_PT(189)
     OR ROM32_INSTR_PT(200) OR ROM32_INSTR_PT(209)
     OR ROM32_INSTR_PT(215) OR ROM32_INSTR_PT(219)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(250)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(259)
     OR ROM32_INSTR_PT(261) OR ROM32_INSTR_PT(262)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(267)
     OR ROM32_INSTR_PT(272) OR ROM32_INSTR_PT(273)
     OR ROM32_INSTR_PT(278) OR ROM32_INSTR_PT(281)
     OR ROM32_INSTR_PT(283) OR ROM32_INSTR_PT(301)
     OR ROM32_INSTR_PT(313) OR ROM32_INSTR_PT(321)
     OR ROM32_INSTR_PT(328) OR ROM32_INSTR_PT(345)
     OR ROM32_INSTR_PT(360) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(368) OR ROM32_INSTR_PT(371)
     OR ROM32_INSTR_PT(390) OR ROM32_INSTR_PT(392)
     OR ROM32_INSTR_PT(396) OR ROM32_INSTR_PT(398)
     OR ROM32_INSTR_PT(401) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(424) OR ROM32_INSTR_PT(433)
     OR ROM32_INSTR_PT(446) OR ROM32_INSTR_PT(468)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(502) OR ROM32_INSTR_PT(519)
     OR ROM32_INSTR_PT(521) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(524) OR ROM32_INSTR_PT(537)
     OR ROM32_INSTR_PT(539) OR ROM32_INSTR_PT(554)
     OR ROM32_INSTR_PT(556) OR ROM32_INSTR_PT(562)
     OR ROM32_INSTR_PT(568) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(583) OR ROM32_INSTR_PT(590)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(595)
     OR ROM32_INSTR_PT(602) OR ROM32_INSTR_PT(607)
     OR ROM32_INSTR_PT(612) OR ROM32_INSTR_PT(614)
     OR ROM32_INSTR_PT(626) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(736)
     OR ROM32_INSTR_PT(762) OR ROM32_INSTR_PT(770)
     OR ROM32_INSTR_PT(870));
MQQ1872:TEMPLATE(17) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(16)
     OR ROM32_INSTR_PT(18) OR ROM32_INSTR_PT(20)
     OR ROM32_INSTR_PT(26) OR ROM32_INSTR_PT(32)
     OR ROM32_INSTR_PT(34) OR ROM32_INSTR_PT(37)
     OR ROM32_INSTR_PT(38) OR ROM32_INSTR_PT(43)
     OR ROM32_INSTR_PT(49) OR ROM32_INSTR_PT(55)
     OR ROM32_INSTR_PT(63) OR ROM32_INSTR_PT(73)
     OR ROM32_INSTR_PT(79) OR ROM32_INSTR_PT(80)
     OR ROM32_INSTR_PT(87) OR ROM32_INSTR_PT(90)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(99)
     OR ROM32_INSTR_PT(103) OR ROM32_INSTR_PT(105)
     OR ROM32_INSTR_PT(112) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(122) OR ROM32_INSTR_PT(127)
     OR ROM32_INSTR_PT(173) OR ROM32_INSTR_PT(184)
     OR ROM32_INSTR_PT(186) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(189) OR ROM32_INSTR_PT(200)
     OR ROM32_INSTR_PT(209) OR ROM32_INSTR_PT(216)
     OR ROM32_INSTR_PT(224) OR ROM32_INSTR_PT(227)
     OR ROM32_INSTR_PT(232) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(250)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(259)
     OR ROM32_INSTR_PT(262) OR ROM32_INSTR_PT(264)
     OR ROM32_INSTR_PT(269) OR ROM32_INSTR_PT(270)
     OR ROM32_INSTR_PT(272) OR ROM32_INSTR_PT(275)
     OR ROM32_INSTR_PT(278) OR ROM32_INSTR_PT(280)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(283)
     OR ROM32_INSTR_PT(284) OR ROM32_INSTR_PT(288)
     OR ROM32_INSTR_PT(299) OR ROM32_INSTR_PT(301)
     OR ROM32_INSTR_PT(303) OR ROM32_INSTR_PT(321)
     OR ROM32_INSTR_PT(326) OR ROM32_INSTR_PT(328)
     OR ROM32_INSTR_PT(340) OR ROM32_INSTR_PT(345)
     OR ROM32_INSTR_PT(348) OR ROM32_INSTR_PT(361)
     OR ROM32_INSTR_PT(366) OR ROM32_INSTR_PT(378)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(383)
     OR ROM32_INSTR_PT(392) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(404)
     OR ROM32_INSTR_PT(406) OR ROM32_INSTR_PT(416)
     OR ROM32_INSTR_PT(418) OR ROM32_INSTR_PT(419)
     OR ROM32_INSTR_PT(421) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(446) OR ROM32_INSTR_PT(468)
     OR ROM32_INSTR_PT(475) OR ROM32_INSTR_PT(476)
     OR ROM32_INSTR_PT(477) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(480)
     OR ROM32_INSTR_PT(481) OR ROM32_INSTR_PT(482)
     OR ROM32_INSTR_PT(490) OR ROM32_INSTR_PT(494)
     OR ROM32_INSTR_PT(497) OR ROM32_INSTR_PT(505)
     OR ROM32_INSTR_PT(508) OR ROM32_INSTR_PT(520)
     OR ROM32_INSTR_PT(521) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(534) OR ROM32_INSTR_PT(535)
     OR ROM32_INSTR_PT(537) OR ROM32_INSTR_PT(538)
     OR ROM32_INSTR_PT(546) OR ROM32_INSTR_PT(547)
     OR ROM32_INSTR_PT(550) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(562)
     OR ROM32_INSTR_PT(574) OR ROM32_INSTR_PT(578)
     OR ROM32_INSTR_PT(582) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(585) OR ROM32_INSTR_PT(591)
     OR ROM32_INSTR_PT(593) OR ROM32_INSTR_PT(598)
     OR ROM32_INSTR_PT(602) OR ROM32_INSTR_PT(606)
     OR ROM32_INSTR_PT(607) OR ROM32_INSTR_PT(608)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(635)
     OR ROM32_INSTR_PT(639) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(647)
     OR ROM32_INSTR_PT(666) OR ROM32_INSTR_PT(677)
     OR ROM32_INSTR_PT(680) OR ROM32_INSTR_PT(698)
     OR ROM32_INSTR_PT(870));
MQQ1873:TEMPLATE(18) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(18)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(34) OR ROM32_INSTR_PT(38)
     OR ROM32_INSTR_PT(49) OR ROM32_INSTR_PT(79)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(111) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(172) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(259)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(396) OR ROM32_INSTR_PT(398)
     OR ROM32_INSTR_PT(424) OR ROM32_INSTR_PT(468)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(537)
     OR ROM32_INSTR_PT(543) OR ROM32_INSTR_PT(554)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(720) OR ROM32_INSTR_PT(807)
     OR ROM32_INSTR_PT(823));
MQQ1874:TEMPLATE(19) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(14)
     OR ROM32_INSTR_PT(18) OR ROM32_INSTR_PT(20)
     OR ROM32_INSTR_PT(23) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(34) OR ROM32_INSTR_PT(38)
     OR ROM32_INSTR_PT(39) OR ROM32_INSTR_PT(42)
     OR ROM32_INSTR_PT(45) OR ROM32_INSTR_PT(49)
     OR ROM32_INSTR_PT(53) OR ROM32_INSTR_PT(57)
     OR ROM32_INSTR_PT(79) OR ROM32_INSTR_PT(85)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(101) OR ROM32_INSTR_PT(102)
     OR ROM32_INSTR_PT(110) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(141) OR ROM32_INSTR_PT(143)
     OR ROM32_INSTR_PT(144) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(178) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(203) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(206) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(232) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(243) OR ROM32_INSTR_PT(251)
     OR ROM32_INSTR_PT(252) OR ROM32_INSTR_PT(258)
     OR ROM32_INSTR_PT(268) OR ROM32_INSTR_PT(271)
     OR ROM32_INSTR_PT(278) OR ROM32_INSTR_PT(281)
     OR ROM32_INSTR_PT(289) OR ROM32_INSTR_PT(294)
     OR ROM32_INSTR_PT(306) OR ROM32_INSTR_PT(323)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(378) OR ROM32_INSTR_PT(382)
     OR ROM32_INSTR_PT(385) OR ROM32_INSTR_PT(386)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(405)
     OR ROM32_INSTR_PT(416) OR ROM32_INSTR_PT(417)
     OR ROM32_INSTR_PT(419) OR ROM32_INSTR_PT(422)
     OR ROM32_INSTR_PT(424) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(435) OR ROM32_INSTR_PT(436)
     OR ROM32_INSTR_PT(452) OR ROM32_INSTR_PT(458)
     OR ROM32_INSTR_PT(468) OR ROM32_INSTR_PT(476)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(507) OR ROM32_INSTR_PT(517)
     OR ROM32_INSTR_PT(521) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(532)
     OR ROM32_INSTR_PT(537) OR ROM32_INSTR_PT(541)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(554)
     OR ROM32_INSTR_PT(569) OR ROM32_INSTR_PT(579)
     OR ROM32_INSTR_PT(581) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(610) OR ROM32_INSTR_PT(615)
     OR ROM32_INSTR_PT(616) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(643) OR ROM32_INSTR_PT(674)
     OR ROM32_INSTR_PT(684) OR ROM32_INSTR_PT(720)
     OR ROM32_INSTR_PT(729) OR ROM32_INSTR_PT(763)
     OR ROM32_INSTR_PT(807) OR ROM32_INSTR_PT(812)
     OR ROM32_INSTR_PT(818) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(823) OR ROM32_INSTR_PT(878)
    );
MQQ1875:TEMPLATE(20) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(12)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(33)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(38)
     OR ROM32_INSTR_PT(42) OR ROM32_INSTR_PT(45)
     OR ROM32_INSTR_PT(49) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(102)
     OR ROM32_INSTR_PT(119) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(196) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(218) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(257)
     OR ROM32_INSTR_PT(258) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(306)
     OR ROM32_INSTR_PT(323) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(362) OR ROM32_INSTR_PT(367)
     OR ROM32_INSTR_PT(382) OR ROM32_INSTR_PT(386)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(396) OR ROM32_INSTR_PT(398)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(422)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(431) OR ROM32_INSTR_PT(435)
     OR ROM32_INSTR_PT(452) OR ROM32_INSTR_PT(454)
     OR ROM32_INSTR_PT(456) OR ROM32_INSTR_PT(464)
     OR ROM32_INSTR_PT(469) OR ROM32_INSTR_PT(472)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(484)
     OR ROM32_INSTR_PT(504) OR ROM32_INSTR_PT(514)
     OR ROM32_INSTR_PT(516) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(537)
     OR ROM32_INSTR_PT(541) OR ROM32_INSTR_PT(543)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(577) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(584) OR ROM32_INSTR_PT(591)
     OR ROM32_INSTR_PT(611) OR ROM32_INSTR_PT(615)
     OR ROM32_INSTR_PT(625) OR ROM32_INSTR_PT(634)
     OR ROM32_INSTR_PT(638) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(684) OR ROM32_INSTR_PT(690)
     OR ROM32_INSTR_PT(718) OR ROM32_INSTR_PT(728)
     OR ROM32_INSTR_PT(751) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(763) OR ROM32_INSTR_PT(805)
     OR ROM32_INSTR_PT(818));
MQQ1876:TEMPLATE(21) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(8) OR ROM32_INSTR_PT(9)
     OR ROM32_INSTR_PT(10) OR ROM32_INSTR_PT(17)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(23)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(38)
     OR ROM32_INSTR_PT(43) OR ROM32_INSTR_PT(60)
     OR ROM32_INSTR_PT(73) OR ROM32_INSTR_PT(74)
     OR ROM32_INSTR_PT(78) OR ROM32_INSTR_PT(80)
     OR ROM32_INSTR_PT(84) OR ROM32_INSTR_PT(87)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(97) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(134) OR ROM32_INSTR_PT(148)
     OR ROM32_INSTR_PT(154) OR ROM32_INSTR_PT(172)
     OR ROM32_INSTR_PT(178) OR ROM32_INSTR_PT(179)
     OR ROM32_INSTR_PT(186) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(194) OR ROM32_INSTR_PT(202)
     OR ROM32_INSTR_PT(206) OR ROM32_INSTR_PT(215)
     OR ROM32_INSTR_PT(218) OR ROM32_INSTR_PT(223)
     OR ROM32_INSTR_PT(224) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(232) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(244) OR ROM32_INSTR_PT(251)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(261)
     OR ROM32_INSTR_PT(262) OR ROM32_INSTR_PT(267)
     OR ROM32_INSTR_PT(270) OR ROM32_INSTR_PT(273)
     OR ROM32_INSTR_PT(275) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(295) OR ROM32_INSTR_PT(297)
     OR ROM32_INSTR_PT(310) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(360)
     OR ROM32_INSTR_PT(362) OR ROM32_INSTR_PT(368)
     OR ROM32_INSTR_PT(371) OR ROM32_INSTR_PT(378)
     OR ROM32_INSTR_PT(385) OR ROM32_INSTR_PT(387)
     OR ROM32_INSTR_PT(390) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(401)
     OR ROM32_INSTR_PT(411) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(416) OR ROM32_INSTR_PT(419)
     OR ROM32_INSTR_PT(421) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(426) OR ROM32_INSTR_PT(433)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(496) OR ROM32_INSTR_PT(502)
     OR ROM32_INSTR_PT(506) OR ROM32_INSTR_PT(507)
     OR ROM32_INSTR_PT(508) OR ROM32_INSTR_PT(516)
     OR ROM32_INSTR_PT(519) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(524) OR ROM32_INSTR_PT(530)
     OR ROM32_INSTR_PT(531) OR ROM32_INSTR_PT(535)
     OR ROM32_INSTR_PT(537) OR ROM32_INSTR_PT(539)
     OR ROM32_INSTR_PT(543) OR ROM32_INSTR_PT(547)
     OR ROM32_INSTR_PT(556) OR ROM32_INSTR_PT(558)
     OR ROM32_INSTR_PT(568) OR ROM32_INSTR_PT(569)
     OR ROM32_INSTR_PT(574) OR ROM32_INSTR_PT(575)
     OR ROM32_INSTR_PT(578) OR ROM32_INSTR_PT(579)
     OR ROM32_INSTR_PT(583) OR ROM32_INSTR_PT(585)
     OR ROM32_INSTR_PT(588) OR ROM32_INSTR_PT(590)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(611)
     OR ROM32_INSTR_PT(612) OR ROM32_INSTR_PT(614)
     OR ROM32_INSTR_PT(621) OR ROM32_INSTR_PT(625)
     OR ROM32_INSTR_PT(626) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(751)
     OR ROM32_INSTR_PT(753) OR ROM32_INSTR_PT(817)
    );
MQQ1877:TEMPLATE(22) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(7)
     OR ROM32_INSTR_PT(8) OR ROM32_INSTR_PT(10)
     OR ROM32_INSTR_PT(12) OR ROM32_INSTR_PT(14)
     OR ROM32_INSTR_PT(17) OR ROM32_INSTR_PT(20)
     OR ROM32_INSTR_PT(23) OR ROM32_INSTR_PT(29)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(38)
     OR ROM32_INSTR_PT(43) OR ROM32_INSTR_PT(53)
     OR ROM32_INSTR_PT(56) OR ROM32_INSTR_PT(57)
     OR ROM32_INSTR_PT(74) OR ROM32_INSTR_PT(78)
     OR ROM32_INSTR_PT(80) OR ROM32_INSTR_PT(93)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(101) OR ROM32_INSTR_PT(114)
     OR ROM32_INSTR_PT(119) OR ROM32_INSTR_PT(122)
     OR ROM32_INSTR_PT(131) OR ROM32_INSTR_PT(134)
     OR ROM32_INSTR_PT(143) OR ROM32_INSTR_PT(148)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(163) OR ROM32_INSTR_PT(164)
     OR ROM32_INSTR_PT(171) OR ROM32_INSTR_PT(172)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(186)
     OR ROM32_INSTR_PT(196) OR ROM32_INSTR_PT(202)
     OR ROM32_INSTR_PT(203) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(207) OR ROM32_INSTR_PT(212)
     OR ROM32_INSTR_PT(218) OR ROM32_INSTR_PT(220)
     OR ROM32_INSTR_PT(223) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(229) OR ROM32_INSTR_PT(243)
     OR ROM32_INSTR_PT(244) OR ROM32_INSTR_PT(251)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(262)
     OR ROM32_INSTR_PT(271) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(295) OR ROM32_INSTR_PT(297)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(310)
     OR ROM32_INSTR_PT(323) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(362) OR ROM32_INSTR_PT(367)
     OR ROM32_INSTR_PT(376) OR ROM32_INSTR_PT(387)
     OR ROM32_INSTR_PT(392) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(396) OR ROM32_INSTR_PT(398)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(411)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(435)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(438)
     OR ROM32_INSTR_PT(452) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(456)
     OR ROM32_INSTR_PT(458) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(464) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(484) OR ROM32_INSTR_PT(486)
     OR ROM32_INSTR_PT(496) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(506) OR ROM32_INSTR_PT(511)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(516)
     OR ROM32_INSTR_PT(517) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(537)
     OR ROM32_INSTR_PT(539) OR ROM32_INSTR_PT(543)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(558)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(575)
     OR ROM32_INSTR_PT(577) OR ROM32_INSTR_PT(580)
     OR ROM32_INSTR_PT(581) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(584) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(601) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(607) OR ROM32_INSTR_PT(611)
     OR ROM32_INSTR_PT(614) OR ROM32_INSTR_PT(622)
     OR ROM32_INSTR_PT(625) OR ROM32_INSTR_PT(634)
     OR ROM32_INSTR_PT(638) OR ROM32_INSTR_PT(643)
     OR ROM32_INSTR_PT(654) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(684) OR ROM32_INSTR_PT(693)
     OR ROM32_INSTR_PT(708) OR ROM32_INSTR_PT(720)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(751)
     OR ROM32_INSTR_PT(753) OR ROM32_INSTR_PT(807)
     OR ROM32_INSTR_PT(817) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(823) OR ROM32_INSTR_PT(845)
     OR ROM32_INSTR_PT(853));
MQQ1878:TEMPLATE(23) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(12) OR ROM32_INSTR_PT(23)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(38)
     OR ROM32_INSTR_PT(56) OR ROM32_INSTR_PT(57)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(111) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(135) OR ROM32_INSTR_PT(143)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(163) OR ROM32_INSTR_PT(179)
     OR ROM32_INSTR_PT(187) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(202) OR ROM32_INSTR_PT(203)
     OR ROM32_INSTR_PT(207) OR ROM32_INSTR_PT(218)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(232) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(243) OR ROM32_INSTR_PT(244)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(254)
     OR ROM32_INSTR_PT(256) OR ROM32_INSTR_PT(257)
     OR ROM32_INSTR_PT(259) OR ROM32_INSTR_PT(260)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(275)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(282)
     OR ROM32_INSTR_PT(293) OR ROM32_INSTR_PT(310)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(362) OR ROM32_INSTR_PT(367)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(378) OR ROM32_INSTR_PT(387)
     OR ROM32_INSTR_PT(394) OR ROM32_INSTR_PT(398)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(416) OR ROM32_INSTR_PT(419)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(434)
     OR ROM32_INSTR_PT(443) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(456)
     OR ROM32_INSTR_PT(458) OR ROM32_INSTR_PT(464)
     OR ROM32_INSTR_PT(469) OR ROM32_INSTR_PT(472)
     OR ROM32_INSTR_PT(484) OR ROM32_INSTR_PT(486)
     OR ROM32_INSTR_PT(501) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(516)
     OR ROM32_INSTR_PT(531) OR ROM32_INSTR_PT(535)
     OR ROM32_INSTR_PT(537) OR ROM32_INSTR_PT(544)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(551)
     OR ROM32_INSTR_PT(557) OR ROM32_INSTR_PT(558)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(577) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(588) OR ROM32_INSTR_PT(591)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(609) OR ROM32_INSTR_PT(611)
     OR ROM32_INSTR_PT(621) OR ROM32_INSTR_PT(625)
     OR ROM32_INSTR_PT(643) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(690) OR ROM32_INSTR_PT(713)
     OR ROM32_INSTR_PT(720) OR ROM32_INSTR_PT(728)
     OR ROM32_INSTR_PT(751) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(807) OR ROM32_INSTR_PT(817)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(823)
     OR ROM32_INSTR_PT(845));
MQQ1879:TEMPLATE(24) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(4)
     OR ROM32_INSTR_PT(5) OR ROM32_INSTR_PT(10)
     OR ROM32_INSTR_PT(13) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(29) OR ROM32_INSTR_PT(34)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(41)
     OR ROM32_INSTR_PT(45) OR ROM32_INSTR_PT(51)
     OR ROM32_INSTR_PT(79) OR ROM32_INSTR_PT(93)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(100)
     OR ROM32_INSTR_PT(106) OR ROM32_INSTR_PT(116)
     OR ROM32_INSTR_PT(124) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(139) OR ROM32_INSTR_PT(142)
     OR ROM32_INSTR_PT(153) OR ROM32_INSTR_PT(159)
     OR ROM32_INSTR_PT(170) OR ROM32_INSTR_PT(172)
     OR ROM32_INSTR_PT(183) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(204) OR ROM32_INSTR_PT(218)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(241) OR ROM32_INSTR_PT(251)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(258)
     OR ROM32_INSTR_PT(260) OR ROM32_INSTR_PT(275)
     OR ROM32_INSTR_PT(276) OR ROM32_INSTR_PT(281)
     OR ROM32_INSTR_PT(282) OR ROM32_INSTR_PT(290)
     OR ROM32_INSTR_PT(293) OR ROM32_INSTR_PT(306)
     OR ROM32_INSTR_PT(309) OR ROM32_INSTR_PT(318)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(362)
     OR ROM32_INSTR_PT(363) OR ROM32_INSTR_PT(374)
     OR ROM32_INSTR_PT(385) OR ROM32_INSTR_PT(393)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(425)
     OR ROM32_INSTR_PT(426) OR ROM32_INSTR_PT(428)
     OR ROM32_INSTR_PT(430) OR ROM32_INSTR_PT(434)
     OR ROM32_INSTR_PT(437) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(454)
     OR ROM32_INSTR_PT(495) OR ROM32_INSTR_PT(501)
     OR ROM32_INSTR_PT(509) OR ROM32_INSTR_PT(516)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(531)
     OR ROM32_INSTR_PT(535) OR ROM32_INSTR_PT(543)
     OR ROM32_INSTR_PT(544) OR ROM32_INSTR_PT(547)
     OR ROM32_INSTR_PT(555) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(574) OR ROM32_INSTR_PT(575)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(587) OR ROM32_INSTR_PT(591)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(609)
     OR ROM32_INSTR_PT(611) OR ROM32_INSTR_PT(615)
     OR ROM32_INSTR_PT(621) OR ROM32_INSTR_PT(624)
     OR ROM32_INSTR_PT(625) OR ROM32_INSTR_PT(646)
     OR ROM32_INSTR_PT(663) OR ROM32_INSTR_PT(690)
     OR ROM32_INSTR_PT(700) OR ROM32_INSTR_PT(729)
     OR ROM32_INSTR_PT(745) OR ROM32_INSTR_PT(763)
     OR ROM32_INSTR_PT(817) OR ROM32_INSTR_PT(845)
    );
MQQ1880:TEMPLATE(25) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(12) OR ROM32_INSTR_PT(20)
     OR ROM32_INSTR_PT(23) OR ROM32_INSTR_PT(35)
     OR ROM32_INSTR_PT(42) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(97) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(119) OR ROM32_INSTR_PT(125)
     OR ROM32_INSTR_PT(132) OR ROM32_INSTR_PT(142)
     OR ROM32_INSTR_PT(143) OR ROM32_INSTR_PT(155)
     OR ROM32_INSTR_PT(158) OR ROM32_INSTR_PT(159)
     OR ROM32_INSTR_PT(163) OR ROM32_INSTR_PT(170)
     OR ROM32_INSTR_PT(172) OR ROM32_INSTR_PT(178)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(194) OR ROM32_INSTR_PT(196)
     OR ROM32_INSTR_PT(203) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(218) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(229) OR ROM32_INSTR_PT(232)
     OR ROM32_INSTR_PT(235) OR ROM32_INSTR_PT(243)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(275)
     OR ROM32_INSTR_PT(276) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(290)
     OR ROM32_INSTR_PT(309) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(362) OR ROM32_INSTR_PT(363)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(378) OR ROM32_INSTR_PT(385)
     OR ROM32_INSTR_PT(394) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(402)
     OR ROM32_INSTR_PT(416) OR ROM32_INSTR_PT(419)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(426) OR ROM32_INSTR_PT(430)
     OR ROM32_INSTR_PT(442) OR ROM32_INSTR_PT(454)
     OR ROM32_INSTR_PT(456) OR ROM32_INSTR_PT(458)
     OR ROM32_INSTR_PT(464) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(474)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(484)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(504) OR ROM32_INSTR_PT(514)
     OR ROM32_INSTR_PT(521) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(531)
     OR ROM32_INSTR_PT(535) OR ROM32_INSTR_PT(541)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(551)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(555)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(575) OR ROM32_INSTR_PT(577)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(611) OR ROM32_INSTR_PT(620)
     OR ROM32_INSTR_PT(629) OR ROM32_INSTR_PT(633)
     OR ROM32_INSTR_PT(642) OR ROM32_INSTR_PT(643)
     OR ROM32_INSTR_PT(654) OR ROM32_INSTR_PT(664)
     OR ROM32_INSTR_PT(690) OR ROM32_INSTR_PT(697)
     OR ROM32_INSTR_PT(708) OR ROM32_INSTR_PT(729)
     OR ROM32_INSTR_PT(731) OR ROM32_INSTR_PT(745)
     OR ROM32_INSTR_PT(792) OR ROM32_INSTR_PT(817)
     OR ROM32_INSTR_PT(818) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(829));
MQQ1881:TEMPLATE(26) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(4)
     OR ROM32_INSTR_PT(5) OR ROM32_INSTR_PT(6)
     OR ROM32_INSTR_PT(8) OR ROM32_INSTR_PT(9)
     OR ROM32_INSTR_PT(10) OR ROM32_INSTR_PT(12)
     OR ROM32_INSTR_PT(13) OR ROM32_INSTR_PT(17)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(23)
     OR ROM32_INSTR_PT(26) OR ROM32_INSTR_PT(29)
     OR ROM32_INSTR_PT(33) OR ROM32_INSTR_PT(35)
     OR ROM32_INSTR_PT(37) OR ROM32_INSTR_PT(39)
     OR ROM32_INSTR_PT(41) OR ROM32_INSTR_PT(43)
     OR ROM32_INSTR_PT(45) OR ROM32_INSTR_PT(49)
     OR ROM32_INSTR_PT(50) OR ROM32_INSTR_PT(51)
     OR ROM32_INSTR_PT(52) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(59)
     OR ROM32_INSTR_PT(60) OR ROM32_INSTR_PT(63)
     OR ROM32_INSTR_PT(66) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(73) OR ROM32_INSTR_PT(74)
     OR ROM32_INSTR_PT(78) OR ROM32_INSTR_PT(80)
     OR ROM32_INSTR_PT(83) OR ROM32_INSTR_PT(84)
     OR ROM32_INSTR_PT(85) OR ROM32_INSTR_PT(87)
     OR ROM32_INSTR_PT(90) OR ROM32_INSTR_PT(92)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(96) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(102) OR ROM32_INSTR_PT(103)
     OR ROM32_INSTR_PT(106) OR ROM32_INSTR_PT(109)
     OR ROM32_INSTR_PT(110) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(124) OR ROM32_INSTR_PT(130)
     OR ROM32_INSTR_PT(134) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(139) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(142) OR ROM32_INSTR_PT(143)
     OR ROM32_INSTR_PT(144) OR ROM32_INSTR_PT(148)
     OR ROM32_INSTR_PT(153) OR ROM32_INSTR_PT(154)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(159) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(169) OR ROM32_INSTR_PT(172)
     OR ROM32_INSTR_PT(174) OR ROM32_INSTR_PT(176)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(180)
     OR ROM32_INSTR_PT(181) OR ROM32_INSTR_PT(183)
     OR ROM32_INSTR_PT(184) OR ROM32_INSTR_PT(186)
     OR ROM32_INSTR_PT(192) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(196) OR ROM32_INSTR_PT(199)
     OR ROM32_INSTR_PT(202) OR ROM32_INSTR_PT(203)
     OR ROM32_INSTR_PT(204) OR ROM32_INSTR_PT(206)
     OR ROM32_INSTR_PT(207) OR ROM32_INSTR_PT(216)
     OR ROM32_INSTR_PT(218) OR ROM32_INSTR_PT(220)
     OR ROM32_INSTR_PT(223) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(233)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(241)
     OR ROM32_INSTR_PT(243) OR ROM32_INSTR_PT(244)
     OR ROM32_INSTR_PT(249) OR ROM32_INSTR_PT(251)
     OR ROM32_INSTR_PT(252) OR ROM32_INSTR_PT(254)
     OR ROM32_INSTR_PT(256) OR ROM32_INSTR_PT(257)
     OR ROM32_INSTR_PT(259) OR ROM32_INSTR_PT(260)
     OR ROM32_INSTR_PT(261) OR ROM32_INSTR_PT(262)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(266)
     OR ROM32_INSTR_PT(267) OR ROM32_INSTR_PT(268)
     OR ROM32_INSTR_PT(269) OR ROM32_INSTR_PT(270)
     OR ROM32_INSTR_PT(273) OR ROM32_INSTR_PT(274)
     OR ROM32_INSTR_PT(275) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(280) OR ROM32_INSTR_PT(281)
     OR ROM32_INSTR_PT(282) OR ROM32_INSTR_PT(284)
     OR ROM32_INSTR_PT(288) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(290) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(306) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(310) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(346)
     OR ROM32_INSTR_PT(348) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(353) OR ROM32_INSTR_PT(356)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(362)
     OR ROM32_INSTR_PT(364) OR ROM32_INSTR_PT(367)
     OR ROM32_INSTR_PT(371) OR ROM32_INSTR_PT(373)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(382) OR ROM32_INSTR_PT(383)
     OR ROM32_INSTR_PT(386) OR ROM32_INSTR_PT(387)
     OR ROM32_INSTR_PT(390) OR ROM32_INSTR_PT(392)
     OR ROM32_INSTR_PT(394) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(400)
     OR ROM32_INSTR_PT(401) OR ROM32_INSTR_PT(402)
     OR ROM32_INSTR_PT(405) OR ROM32_INSTR_PT(406)
     OR ROM32_INSTR_PT(409) OR ROM32_INSTR_PT(411)
     OR ROM32_INSTR_PT(412) OR ROM32_INSTR_PT(415)
     OR ROM32_INSTR_PT(417) OR ROM32_INSTR_PT(421)
     OR ROM32_INSTR_PT(422) OR ROM32_INSTR_PT(423)
     OR ROM32_INSTR_PT(424) OR ROM32_INSTR_PT(425)
     OR ROM32_INSTR_PT(426) OR ROM32_INSTR_PT(428)
     OR ROM32_INSTR_PT(431) OR ROM32_INSTR_PT(433)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(437)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(458)
     OR ROM32_INSTR_PT(459) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(464) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(475)
     OR ROM32_INSTR_PT(478) OR ROM32_INSTR_PT(479)
     OR ROM32_INSTR_PT(481) OR ROM32_INSTR_PT(482)
     OR ROM32_INSTR_PT(484) OR ROM32_INSTR_PT(486)
     OR ROM32_INSTR_PT(490) OR ROM32_INSTR_PT(491)
     OR ROM32_INSTR_PT(494) OR ROM32_INSTR_PT(495)
     OR ROM32_INSTR_PT(496) OR ROM32_INSTR_PT(501)
     OR ROM32_INSTR_PT(502) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(506) OR ROM32_INSTR_PT(507)
     OR ROM32_INSTR_PT(508) OR ROM32_INSTR_PT(509)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(516)
     OR ROM32_INSTR_PT(519) OR ROM32_INSTR_PT(520)
     OR ROM32_INSTR_PT(521) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(524) OR ROM32_INSTR_PT(530)
     OR ROM32_INSTR_PT(531) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(535) OR ROM32_INSTR_PT(539)
     OR ROM32_INSTR_PT(543) OR ROM32_INSTR_PT(544)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(550)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(555)
     OR ROM32_INSTR_PT(556) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(568) OR ROM32_INSTR_PT(569)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(575) OR ROM32_INSTR_PT(578)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(582) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(585) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(590) OR ROM32_INSTR_PT(591)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(602)
     OR ROM32_INSTR_PT(603) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(609) OR ROM32_INSTR_PT(610)
     OR ROM32_INSTR_PT(611) OR ROM32_INSTR_PT(612)
     OR ROM32_INSTR_PT(613) OR ROM32_INSTR_PT(614)
     OR ROM32_INSTR_PT(615) OR ROM32_INSTR_PT(621)
     OR ROM32_INSTR_PT(624) OR ROM32_INSTR_PT(625)
     OR ROM32_INSTR_PT(626) OR ROM32_INSTR_PT(629)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(639)
     OR ROM32_INSTR_PT(640) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(643) OR ROM32_INSTR_PT(654)
     OR ROM32_INSTR_PT(660) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(664) OR ROM32_INSTR_PT(666)
     OR ROM32_INSTR_PT(674) OR ROM32_INSTR_PT(677)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(697)
     OR ROM32_INSTR_PT(708) OR ROM32_INSTR_PT(711)
     OR ROM32_INSTR_PT(713) OR ROM32_INSTR_PT(718)
     OR ROM32_INSTR_PT(719) OR ROM32_INSTR_PT(720)
     OR ROM32_INSTR_PT(729) OR ROM32_INSTR_PT(755)
     OR ROM32_INSTR_PT(763) OR ROM32_INSTR_PT(792)
     OR ROM32_INSTR_PT(805) OR ROM32_INSTR_PT(807)
     OR ROM32_INSTR_PT(812) OR ROM32_INSTR_PT(817)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(823)
     OR ROM32_INSTR_PT(829) OR ROM32_INSTR_PT(831)
     OR ROM32_INSTR_PT(845) OR ROM32_INSTR_PT(854)
     OR ROM32_INSTR_PT(855) OR ROM32_INSTR_PT(857)
     OR ROM32_INSTR_PT(862) OR ROM32_INSTR_PT(870)
     OR ROM32_INSTR_PT(872) OR ROM32_INSTR_PT(878)
    );
MQQ1882:TEMPLATE(27) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(7)
     OR ROM32_INSTR_PT(8) OR ROM32_INSTR_PT(9)
     OR ROM32_INSTR_PT(10) OR ROM32_INSTR_PT(12)
     OR ROM32_INSTR_PT(14) OR ROM32_INSTR_PT(17)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(33) OR ROM32_INSTR_PT(37)
     OR ROM32_INSTR_PT(39) OR ROM32_INSTR_PT(42)
     OR ROM32_INSTR_PT(45) OR ROM32_INSTR_PT(49)
     OR ROM32_INSTR_PT(52) OR ROM32_INSTR_PT(53)
     OR ROM32_INSTR_PT(56) OR ROM32_INSTR_PT(57)
     OR ROM32_INSTR_PT(59) OR ROM32_INSTR_PT(63)
     OR ROM32_INSTR_PT(66) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(74) OR ROM32_INSTR_PT(83)
     OR ROM32_INSTR_PT(84) OR ROM32_INSTR_PT(85)
     OR ROM32_INSTR_PT(90) OR ROM32_INSTR_PT(93)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(96)
     OR ROM32_INSTR_PT(101) OR ROM32_INSTR_PT(102)
     OR ROM32_INSTR_PT(103) OR ROM32_INSTR_PT(109)
     OR ROM32_INSTR_PT(110) OR ROM32_INSTR_PT(114)
     OR ROM32_INSTR_PT(115) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(130) OR ROM32_INSTR_PT(131)
     OR ROM32_INSTR_PT(134) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(142) OR ROM32_INSTR_PT(143)
     OR ROM32_INSTR_PT(144) OR ROM32_INSTR_PT(148)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(159) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(164) OR ROM32_INSTR_PT(169)
     OR ROM32_INSTR_PT(170) OR ROM32_INSTR_PT(171)
     OR ROM32_INSTR_PT(176) OR ROM32_INSTR_PT(178)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(180)
     OR ROM32_INSTR_PT(181) OR ROM32_INSTR_PT(184)
     OR ROM32_INSTR_PT(187) OR ROM32_INSTR_PT(192)
     OR ROM32_INSTR_PT(194) OR ROM32_INSTR_PT(196)
     OR ROM32_INSTR_PT(199) OR ROM32_INSTR_PT(202)
     OR ROM32_INSTR_PT(203) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(206) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(212) OR ROM32_INSTR_PT(216)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(223)
     OR ROM32_INSTR_PT(224) OR ROM32_INSTR_PT(227)
     OR ROM32_INSTR_PT(232) OR ROM32_INSTR_PT(233)
     OR ROM32_INSTR_PT(235) OR ROM32_INSTR_PT(238)
     OR ROM32_INSTR_PT(240) OR ROM32_INSTR_PT(243)
     OR ROM32_INSTR_PT(244) OR ROM32_INSTR_PT(249)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(252)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(259) OR ROM32_INSTR_PT(261)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(266)
     OR ROM32_INSTR_PT(267) OR ROM32_INSTR_PT(268)
     OR ROM32_INSTR_PT(269) OR ROM32_INSTR_PT(271)
     OR ROM32_INSTR_PT(274) OR ROM32_INSTR_PT(276)
     OR ROM32_INSTR_PT(278) OR ROM32_INSTR_PT(280)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(284)
     OR ROM32_INSTR_PT(288) OR ROM32_INSTR_PT(290)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(310) OR ROM32_INSTR_PT(323)
     OR ROM32_INSTR_PT(335) OR ROM32_INSTR_PT(344)
     OR ROM32_INSTR_PT(348) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(363)
     OR ROM32_INSTR_PT(364) OR ROM32_INSTR_PT(367)
     OR ROM32_INSTR_PT(371) OR ROM32_INSTR_PT(373)
     OR ROM32_INSTR_PT(376) OR ROM32_INSTR_PT(378)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(382) OR ROM32_INSTR_PT(383)
     OR ROM32_INSTR_PT(386) OR ROM32_INSTR_PT(390)
     OR ROM32_INSTR_PT(392) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(395) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(400)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(405)
     OR ROM32_INSTR_PT(406) OR ROM32_INSTR_PT(411)
     OR ROM32_INSTR_PT(416) OR ROM32_INSTR_PT(417)
     OR ROM32_INSTR_PT(419) OR ROM32_INSTR_PT(422)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(425) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(430) OR ROM32_INSTR_PT(431)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(435)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(438)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(442)
     OR ROM32_INSTR_PT(452) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(456) OR ROM32_INSTR_PT(458)
     OR ROM32_INSTR_PT(464) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(474)
     OR ROM32_INSTR_PT(475) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(481)
     OR ROM32_INSTR_PT(482) OR ROM32_INSTR_PT(484)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(494)
     OR ROM32_INSTR_PT(503) OR ROM32_INSTR_PT(506)
     OR ROM32_INSTR_PT(507) OR ROM32_INSTR_PT(511)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(517)
     OR ROM32_INSTR_PT(520) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(524)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(531)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(541) OR ROM32_INSTR_PT(550)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(555)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(569)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(575)
     OR ROM32_INSTR_PT(577) OR ROM32_INSTR_PT(579)
     OR ROM32_INSTR_PT(580) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(582) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(584) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(601) OR ROM32_INSTR_PT(602)
     OR ROM32_INSTR_PT(605) OR ROM32_INSTR_PT(610)
     OR ROM32_INSTR_PT(615) OR ROM32_INSTR_PT(620)
     OR ROM32_INSTR_PT(622) OR ROM32_INSTR_PT(626)
     OR ROM32_INSTR_PT(629) OR ROM32_INSTR_PT(630)
     OR ROM32_INSTR_PT(634) OR ROM32_INSTR_PT(638)
     OR ROM32_INSTR_PT(639) OR ROM32_INSTR_PT(640)
     OR ROM32_INSTR_PT(642) OR ROM32_INSTR_PT(643)
     OR ROM32_INSTR_PT(654) OR ROM32_INSTR_PT(660)
     OR ROM32_INSTR_PT(663) OR ROM32_INSTR_PT(664)
     OR ROM32_INSTR_PT(666) OR ROM32_INSTR_PT(674)
     OR ROM32_INSTR_PT(677) OR ROM32_INSTR_PT(684)
     OR ROM32_INSTR_PT(693) OR ROM32_INSTR_PT(697)
     OR ROM32_INSTR_PT(708) OR ROM32_INSTR_PT(719)
     OR ROM32_INSTR_PT(720) OR ROM32_INSTR_PT(729)
     OR ROM32_INSTR_PT(745) OR ROM32_INSTR_PT(755)
     OR ROM32_INSTR_PT(763) OR ROM32_INSTR_PT(792)
     OR ROM32_INSTR_PT(805) OR ROM32_INSTR_PT(807)
     OR ROM32_INSTR_PT(812) OR ROM32_INSTR_PT(818)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(823)
     OR ROM32_INSTR_PT(829) OR ROM32_INSTR_PT(831)
     OR ROM32_INSTR_PT(853) OR ROM32_INSTR_PT(854)
     OR ROM32_INSTR_PT(855) OR ROM32_INSTR_PT(862)
     OR ROM32_INSTR_PT(870) OR ROM32_INSTR_PT(878)
    );
MQQ1883:TEMPLATE(28) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(4)
     OR ROM32_INSTR_PT(5) OR ROM32_INSTR_PT(8)
     OR ROM32_INSTR_PT(9) OR ROM32_INSTR_PT(12)
     OR ROM32_INSTR_PT(13) OR ROM32_INSTR_PT(16)
     OR ROM32_INSTR_PT(17) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(32) OR ROM32_INSTR_PT(37)
     OR ROM32_INSTR_PT(39) OR ROM32_INSTR_PT(41)
     OR ROM32_INSTR_PT(45) OR ROM32_INSTR_PT(51)
     OR ROM32_INSTR_PT(52) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(59)
     OR ROM32_INSTR_PT(63) OR ROM32_INSTR_PT(66)
     OR ROM32_INSTR_PT(67) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(73) OR ROM32_INSTR_PT(74)
     OR ROM32_INSTR_PT(77) OR ROM32_INSTR_PT(83)
     OR ROM32_INSTR_PT(84) OR ROM32_INSTR_PT(85)
     OR ROM32_INSTR_PT(87) OR ROM32_INSTR_PT(90)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(98) OR ROM32_INSTR_PT(99)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(102) OR ROM32_INSTR_PT(103)
     OR ROM32_INSTR_PT(106) OR ROM32_INSTR_PT(109)
     OR ROM32_INSTR_PT(114) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(118)
     OR ROM32_INSTR_PT(124) OR ROM32_INSTR_PT(125)
     OR ROM32_INSTR_PT(127) OR ROM32_INSTR_PT(132)
     OR ROM32_INSTR_PT(134) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(139) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(142) OR ROM32_INSTR_PT(143)
     OR ROM32_INSTR_PT(148) OR ROM32_INSTR_PT(153)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(159) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(169) OR ROM32_INSTR_PT(171)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(183)
     OR ROM32_INSTR_PT(184) OR ROM32_INSTR_PT(192)
     OR ROM32_INSTR_PT(194) OR ROM32_INSTR_PT(196)
     OR ROM32_INSTR_PT(199) OR ROM32_INSTR_PT(200)
     OR ROM32_INSTR_PT(202) OR ROM32_INSTR_PT(203)
     OR ROM32_INSTR_PT(204) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(216) OR ROM32_INSTR_PT(219)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(223)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(238)
     OR ROM32_INSTR_PT(241) OR ROM32_INSTR_PT(243)
     OR ROM32_INSTR_PT(249) OR ROM32_INSTR_PT(250)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(254)
     OR ROM32_INSTR_PT(256) OR ROM32_INSTR_PT(259)
     OR ROM32_INSTR_PT(260) OR ROM32_INSTR_PT(261)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(266)
     OR ROM32_INSTR_PT(267) OR ROM32_INSTR_PT(268)
     OR ROM32_INSTR_PT(269) OR ROM32_INSTR_PT(270)
     OR ROM32_INSTR_PT(273) OR ROM32_INSTR_PT(280)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(282)
     OR ROM32_INSTR_PT(284) OR ROM32_INSTR_PT(288)
     OR ROM32_INSTR_PT(290) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(306) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(313) OR ROM32_INSTR_PT(318)
     OR ROM32_INSTR_PT(328) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(348)
     OR ROM32_INSTR_PT(350) OR ROM32_INSTR_PT(361)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(371)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(382) OR ROM32_INSTR_PT(383)
     OR ROM32_INSTR_PT(386) OR ROM32_INSTR_PT(390)
     OR ROM32_INSTR_PT(392) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(401)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(406)
     OR ROM32_INSTR_PT(409) OR ROM32_INSTR_PT(411)
     OR ROM32_INSTR_PT(412) OR ROM32_INSTR_PT(415)
     OR ROM32_INSTR_PT(421) OR ROM32_INSTR_PT(422)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(425)
     OR ROM32_INSTR_PT(426) OR ROM32_INSTR_PT(428)
     OR ROM32_INSTR_PT(431) OR ROM32_INSTR_PT(433)
     OR ROM32_INSTR_PT(437) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(458) OR ROM32_INSTR_PT(464)
     OR ROM32_INSTR_PT(469) OR ROM32_INSTR_PT(472)
     OR ROM32_INSTR_PT(475) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(481)
     OR ROM32_INSTR_PT(482) OR ROM32_INSTR_PT(484)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(491) OR ROM32_INSTR_PT(494)
     OR ROM32_INSTR_PT(495) OR ROM32_INSTR_PT(501)
     OR ROM32_INSTR_PT(502) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(504) OR ROM32_INSTR_PT(506)
     OR ROM32_INSTR_PT(508) OR ROM32_INSTR_PT(509)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(519)
     OR ROM32_INSTR_PT(520) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(524) OR ROM32_INSTR_PT(530)
     OR ROM32_INSTR_PT(531) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(544) OR ROM32_INSTR_PT(550)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(555)
     OR ROM32_INSTR_PT(556) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(568) OR ROM32_INSTR_PT(578)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(582) OR ROM32_INSTR_PT(585)
     OR ROM32_INSTR_PT(588) OR ROM32_INSTR_PT(590)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(595)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(602)
     OR ROM32_INSTR_PT(605) OR ROM32_INSTR_PT(609)
     OR ROM32_INSTR_PT(612) OR ROM32_INSTR_PT(613)
     OR ROM32_INSTR_PT(615) OR ROM32_INSTR_PT(621)
     OR ROM32_INSTR_PT(624) OR ROM32_INSTR_PT(626)
     OR ROM32_INSTR_PT(629) OR ROM32_INSTR_PT(630)
     OR ROM32_INSTR_PT(639) OR ROM32_INSTR_PT(640)
     OR ROM32_INSTR_PT(642) OR ROM32_INSTR_PT(643)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(654)
     OR ROM32_INSTR_PT(660) OR ROM32_INSTR_PT(664)
     OR ROM32_INSTR_PT(666) OR ROM32_INSTR_PT(674)
     OR ROM32_INSTR_PT(677) OR ROM32_INSTR_PT(697)
     OR ROM32_INSTR_PT(708) OR ROM32_INSTR_PT(719)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(729)
     OR ROM32_INSTR_PT(731) OR ROM32_INSTR_PT(736)
     OR ROM32_INSTR_PT(751) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(755) OR ROM32_INSTR_PT(762)
     OR ROM32_INSTR_PT(763) OR ROM32_INSTR_PT(770)
     OR ROM32_INSTR_PT(792) OR ROM32_INSTR_PT(805)
     OR ROM32_INSTR_PT(812) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(829) OR ROM32_INSTR_PT(854)
     OR ROM32_INSTR_PT(855) OR ROM32_INSTR_PT(862)
     OR ROM32_INSTR_PT(870) OR ROM32_INSTR_PT(878)
    );
MQQ1884:TEMPLATE(29) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(4)
     OR ROM32_INSTR_PT(5) OR ROM32_INSTR_PT(6)
     OR ROM32_INSTR_PT(7) OR ROM32_INSTR_PT(8)
     OR ROM32_INSTR_PT(9) OR ROM32_INSTR_PT(10)
     OR ROM32_INSTR_PT(13) OR ROM32_INSTR_PT(14)
     OR ROM32_INSTR_PT(16) OR ROM32_INSTR_PT(17)
     OR ROM32_INSTR_PT(23) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(27) OR ROM32_INSTR_PT(30)
     OR ROM32_INSTR_PT(37) OR ROM32_INSTR_PT(41)
     OR ROM32_INSTR_PT(49) OR ROM32_INSTR_PT(51)
     OR ROM32_INSTR_PT(52) OR ROM32_INSTR_PT(53)
     OR ROM32_INSTR_PT(59) OR ROM32_INSTR_PT(63)
     OR ROM32_INSTR_PT(66) OR ROM32_INSTR_PT(67)
     OR ROM32_INSTR_PT(73) OR ROM32_INSTR_PT(74)
     OR ROM32_INSTR_PT(77) OR ROM32_INSTR_PT(78)
     OR ROM32_INSTR_PT(84) OR ROM32_INSTR_PT(87)
     OR ROM32_INSTR_PT(90) OR ROM32_INSTR_PT(93)
     OR ROM32_INSTR_PT(97) OR ROM32_INSTR_PT(99)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(103)
     OR ROM32_INSTR_PT(106) OR ROM32_INSTR_PT(114)
     OR ROM32_INSTR_PT(115) OR ROM32_INSTR_PT(116)
     OR ROM32_INSTR_PT(117) OR ROM32_INSTR_PT(118)
     OR ROM32_INSTR_PT(124) OR ROM32_INSTR_PT(127)
     OR ROM32_INSTR_PT(130) OR ROM32_INSTR_PT(131)
     OR ROM32_INSTR_PT(132) OR ROM32_INSTR_PT(134)
     OR ROM32_INSTR_PT(135) OR ROM32_INSTR_PT(139)
     OR ROM32_INSTR_PT(148) OR ROM32_INSTR_PT(153)
     OR ROM32_INSTR_PT(159) OR ROM32_INSTR_PT(164)
     OR ROM32_INSTR_PT(169) OR ROM32_INSTR_PT(171)
     OR ROM32_INSTR_PT(172) OR ROM32_INSTR_PT(181)
     OR ROM32_INSTR_PT(183) OR ROM32_INSTR_PT(184)
     OR ROM32_INSTR_PT(187) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(200) OR ROM32_INSTR_PT(204)
     OR ROM32_INSTR_PT(205) OR ROM32_INSTR_PT(212)
     OR ROM32_INSTR_PT(216) OR ROM32_INSTR_PT(219)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(223)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(232) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(241)
     OR ROM32_INSTR_PT(244) OR ROM32_INSTR_PT(250)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(259) OR ROM32_INSTR_PT(260)
     OR ROM32_INSTR_PT(261) OR ROM32_INSTR_PT(264)
     OR ROM32_INSTR_PT(267) OR ROM32_INSTR_PT(269)
     OR ROM32_INSTR_PT(270) OR ROM32_INSTR_PT(271)
     OR ROM32_INSTR_PT(273) OR ROM32_INSTR_PT(274)
     OR ROM32_INSTR_PT(275) OR ROM32_INSTR_PT(280)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(282)
     OR ROM32_INSTR_PT(284) OR ROM32_INSTR_PT(288)
     OR ROM32_INSTR_PT(289) OR ROM32_INSTR_PT(290)
     OR ROM32_INSTR_PT(293) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(306) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(310) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(322)
     OR ROM32_INSTR_PT(323) OR ROM32_INSTR_PT(328)
     OR ROM32_INSTR_PT(337) OR ROM32_INSTR_PT(348)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(371)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(378)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(383) OR ROM32_INSTR_PT(387)
     OR ROM32_INSTR_PT(390) OR ROM32_INSTR_PT(392)
     OR ROM32_INSTR_PT(393) OR ROM32_INSTR_PT(398)
     OR ROM32_INSTR_PT(400) OR ROM32_INSTR_PT(401)
     OR ROM32_INSTR_PT(406) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(411) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(416)
     OR ROM32_INSTR_PT(419) OR ROM32_INSTR_PT(421)
     OR ROM32_INSTR_PT(425) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(428) OR ROM32_INSTR_PT(433)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(435)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(437)
     OR ROM32_INSTR_PT(438) OR ROM32_INSTR_PT(441)
     OR ROM32_INSTR_PT(443) OR ROM32_INSTR_PT(451)
     OR ROM32_INSTR_PT(452) OR ROM32_INSTR_PT(465)
     OR ROM32_INSTR_PT(475) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(481)
     OR ROM32_INSTR_PT(482) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(494) OR ROM32_INSTR_PT(495)
     OR ROM32_INSTR_PT(501) OR ROM32_INSTR_PT(502)
     OR ROM32_INSTR_PT(506) OR ROM32_INSTR_PT(507)
     OR ROM32_INSTR_PT(508) OR ROM32_INSTR_PT(509)
     OR ROM32_INSTR_PT(511) OR ROM32_INSTR_PT(517)
     OR ROM32_INSTR_PT(519) OR ROM32_INSTR_PT(520)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(524)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(531)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(535) OR ROM32_INSTR_PT(543)
     OR ROM32_INSTR_PT(544) OR ROM32_INSTR_PT(547)
     OR ROM32_INSTR_PT(550) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(556)
     OR ROM32_INSTR_PT(557) OR ROM32_INSTR_PT(558)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(568)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(575) OR ROM32_INSTR_PT(578)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(580)
     OR ROM32_INSTR_PT(581) OR ROM32_INSTR_PT(582)
     OR ROM32_INSTR_PT(584) OR ROM32_INSTR_PT(585)
     OR ROM32_INSTR_PT(587) OR ROM32_INSTR_PT(590)
     OR ROM32_INSTR_PT(595) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(601)
     OR ROM32_INSTR_PT(602) OR ROM32_INSTR_PT(609)
     OR ROM32_INSTR_PT(612) OR ROM32_INSTR_PT(622)
     OR ROM32_INSTR_PT(624) OR ROM32_INSTR_PT(625)
     OR ROM32_INSTR_PT(626) OR ROM32_INSTR_PT(629)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(634)
     OR ROM32_INSTR_PT(638) OR ROM32_INSTR_PT(639)
     OR ROM32_INSTR_PT(640) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(664) OR ROM32_INSTR_PT(666)
     OR ROM32_INSTR_PT(677) OR ROM32_INSTR_PT(684)
     OR ROM32_INSTR_PT(693) OR ROM32_INSTR_PT(697)
     OR ROM32_INSTR_PT(719) OR ROM32_INSTR_PT(726)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(736)
     OR ROM32_INSTR_PT(751) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(755) OR ROM32_INSTR_PT(762)
     OR ROM32_INSTR_PT(770) OR ROM32_INSTR_PT(792)
     OR ROM32_INSTR_PT(829) OR ROM32_INSTR_PT(845)
     OR ROM32_INSTR_PT(853) OR ROM32_INSTR_PT(855)
     OR ROM32_INSTR_PT(862) OR ROM32_INSTR_PT(870)
    );
MQQ1885:TEMPLATE(30) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(4)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(8)
     OR ROM32_INSTR_PT(9) OR ROM32_INSTR_PT(13)
     OR ROM32_INSTR_PT(16) OR ROM32_INSTR_PT(17)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(32) OR ROM32_INSTR_PT(37)
     OR ROM32_INSTR_PT(41) OR ROM32_INSTR_PT(45)
     OR ROM32_INSTR_PT(49) OR ROM32_INSTR_PT(50)
     OR ROM32_INSTR_PT(51) OR ROM32_INSTR_PT(52)
     OR ROM32_INSTR_PT(55) OR ROM32_INSTR_PT(59)
     OR ROM32_INSTR_PT(63) OR ROM32_INSTR_PT(66)
     OR ROM32_INSTR_PT(67) OR ROM32_INSTR_PT(73)
     OR ROM32_INSTR_PT(74) OR ROM32_INSTR_PT(77)
     OR ROM32_INSTR_PT(78) OR ROM32_INSTR_PT(79)
     OR ROM32_INSTR_PT(80) OR ROM32_INSTR_PT(84)
     OR ROM32_INSTR_PT(85) OR ROM32_INSTR_PT(87)
     OR ROM32_INSTR_PT(90) OR ROM32_INSTR_PT(92)
     OR ROM32_INSTR_PT(99) OR ROM32_INSTR_PT(100)
     OR ROM32_INSTR_PT(103) OR ROM32_INSTR_PT(105)
     OR ROM32_INSTR_PT(106) OR ROM32_INSTR_PT(111)
     OR ROM32_INSTR_PT(114) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(122) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(127) OR ROM32_INSTR_PT(130)
     OR ROM32_INSTR_PT(134) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(139) OR ROM32_INSTR_PT(142)
     OR ROM32_INSTR_PT(148) OR ROM32_INSTR_PT(153)
     OR ROM32_INSTR_PT(169) OR ROM32_INSTR_PT(171)
     OR ROM32_INSTR_PT(176) OR ROM32_INSTR_PT(179)
     OR ROM32_INSTR_PT(180) OR ROM32_INSTR_PT(181)
     OR ROM32_INSTR_PT(183) OR ROM32_INSTR_PT(184)
     OR ROM32_INSTR_PT(186) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(200) OR ROM32_INSTR_PT(204)
     OR ROM32_INSTR_PT(209) OR ROM32_INSTR_PT(214)
     OR ROM32_INSTR_PT(215) OR ROM32_INSTR_PT(216)
     OR ROM32_INSTR_PT(219) OR ROM32_INSTR_PT(220)
     OR ROM32_INSTR_PT(222) OR ROM32_INSTR_PT(223)
     OR ROM32_INSTR_PT(224) OR ROM32_INSTR_PT(227)
     OR ROM32_INSTR_PT(229) OR ROM32_INSTR_PT(233)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(241)
     OR ROM32_INSTR_PT(250) OR ROM32_INSTR_PT(254)
     OR ROM32_INSTR_PT(256) OR ROM32_INSTR_PT(259)
     OR ROM32_INSTR_PT(260) OR ROM32_INSTR_PT(261)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(267)
     OR ROM32_INSTR_PT(269) OR ROM32_INSTR_PT(270)
     OR ROM32_INSTR_PT(272) OR ROM32_INSTR_PT(273)
     OR ROM32_INSTR_PT(274) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(280) OR ROM32_INSTR_PT(282)
     OR ROM32_INSTR_PT(283) OR ROM32_INSTR_PT(288)
     OR ROM32_INSTR_PT(293) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(306) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(321)
     OR ROM32_INSTR_PT(328) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(343) OR ROM32_INSTR_PT(345)
     OR ROM32_INSTR_PT(346) OR ROM32_INSTR_PT(348)
     OR ROM32_INSTR_PT(356) OR ROM32_INSTR_PT(361)
     OR ROM32_INSTR_PT(364) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(368) OR ROM32_INSTR_PT(371)
     OR ROM32_INSTR_PT(373) OR ROM32_INSTR_PT(374)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(383)
     OR ROM32_INSTR_PT(390) OR ROM32_INSTR_PT(392)
     OR ROM32_INSTR_PT(393) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(400) OR ROM32_INSTR_PT(401)
     OR ROM32_INSTR_PT(406) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(411) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(421)
     OR ROM32_INSTR_PT(424) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(428) OR ROM32_INSTR_PT(431)
     OR ROM32_INSTR_PT(433) OR ROM32_INSTR_PT(437)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(459)
     OR ROM32_INSTR_PT(461) OR ROM32_INSTR_PT(475)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(481)
     OR ROM32_INSTR_PT(482) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(494) OR ROM32_INSTR_PT(495)
     OR ROM32_INSTR_PT(501) OR ROM32_INSTR_PT(502)
     OR ROM32_INSTR_PT(506) OR ROM32_INSTR_PT(507)
     OR ROM32_INSTR_PT(508) OR ROM32_INSTR_PT(509)
     OR ROM32_INSTR_PT(519) OR ROM32_INSTR_PT(520)
     OR ROM32_INSTR_PT(521) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(524) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(539) OR ROM32_INSTR_PT(544)
     OR ROM32_INSTR_PT(550) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(555)
     OR ROM32_INSTR_PT(556) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(562)
     OR ROM32_INSTR_PT(568) OR ROM32_INSTR_PT(570)
     OR ROM32_INSTR_PT(575) OR ROM32_INSTR_PT(578)
     OR ROM32_INSTR_PT(581) OR ROM32_INSTR_PT(582)
     OR ROM32_INSTR_PT(583) OR ROM32_INSTR_PT(585)
     OR ROM32_INSTR_PT(587) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(590) OR ROM32_INSTR_PT(595)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(602)
     OR ROM32_INSTR_PT(603) OR ROM32_INSTR_PT(607)
     OR ROM32_INSTR_PT(609) OR ROM32_INSTR_PT(612)
     OR ROM32_INSTR_PT(615) OR ROM32_INSTR_PT(624)
     OR ROM32_INSTR_PT(626) OR ROM32_INSTR_PT(629)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(639)
     OR ROM32_INSTR_PT(640) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(666)
     OR ROM32_INSTR_PT(677) OR ROM32_INSTR_PT(683)
     OR ROM32_INSTR_PT(685) OR ROM32_INSTR_PT(689)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(711)
     OR ROM32_INSTR_PT(719) OR ROM32_INSTR_PT(720)
     OR ROM32_INSTR_PT(726) OR ROM32_INSTR_PT(728)
     OR ROM32_INSTR_PT(729) OR ROM32_INSTR_PT(736)
     OR ROM32_INSTR_PT(751) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(755) OR ROM32_INSTR_PT(762)
     OR ROM32_INSTR_PT(763) OR ROM32_INSTR_PT(770)
     OR ROM32_INSTR_PT(807) OR ROM32_INSTR_PT(823)
     OR ROM32_INSTR_PT(831) OR ROM32_INSTR_PT(845)
     OR ROM32_INSTR_PT(855) OR ROM32_INSTR_PT(862)
     OR ROM32_INSTR_PT(870));
MQQ1886:TEMPLATE(31) <= 
    (ROM32_INSTR_PT(31) OR ROM32_INSTR_PT(62)
     OR ROM32_INSTR_PT(81) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(104) OR ROM32_INSTR_PT(145)
     OR ROM32_INSTR_PT(147) OR ROM32_INSTR_PT(150)
     OR ROM32_INSTR_PT(162) OR ROM32_INSTR_PT(175)
     OR ROM32_INSTR_PT(185) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(208) OR ROM32_INSTR_PT(210)
     OR ROM32_INSTR_PT(225) OR ROM32_INSTR_PT(228)
     OR ROM32_INSTR_PT(230) OR ROM32_INSTR_PT(232)
     OR ROM32_INSTR_PT(235) OR ROM32_INSTR_PT(245)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(279)
     OR ROM32_INSTR_PT(285) OR ROM32_INSTR_PT(292)
     OR ROM32_INSTR_PT(302) OR ROM32_INSTR_PT(307)
     OR ROM32_INSTR_PT(312) OR ROM32_INSTR_PT(325)
     OR ROM32_INSTR_PT(329) OR ROM32_INSTR_PT(338)
     OR ROM32_INSTR_PT(378) OR ROM32_INSTR_PT(398)
     OR ROM32_INSTR_PT(416) OR ROM32_INSTR_PT(419)
     OR ROM32_INSTR_PT(463) OR ROM32_INSTR_PT(489)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(629)
     OR ROM32_INSTR_PT(632) OR ROM32_INSTR_PT(640)
     OR ROM32_INSTR_PT(641) OR ROM32_INSTR_PT(653)
     OR ROM32_INSTR_PT(672) OR ROM32_INSTR_PT(720)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(751)
     OR ROM32_INSTR_PT(752) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(759) OR ROM32_INSTR_PT(774)
     OR ROM32_INSTR_PT(787) OR ROM32_INSTR_PT(803)
     OR ROM32_INSTR_PT(807) OR ROM32_INSTR_PT(823)
    );
MQQ1887:UCODE_END <= 
    (ROM32_INSTR_PT(198) OR ROM32_INSTR_PT(201)
     OR ROM32_INSTR_PT(213) OR ROM32_INSTR_PT(384)
     OR ROM32_INSTR_PT(438) OR ROM32_INSTR_PT(440)
     OR ROM32_INSTR_PT(450) OR ROM32_INSTR_PT(513)
     OR ROM32_INSTR_PT(515) OR ROM32_INSTR_PT(528)
     OR ROM32_INSTR_PT(541) OR ROM32_INSTR_PT(548)
     OR ROM32_INSTR_PT(553) OR ROM32_INSTR_PT(559)
     OR ROM32_INSTR_PT(567) OR ROM32_INSTR_PT(573)
     OR ROM32_INSTR_PT(576) OR ROM32_INSTR_PT(580)
     OR ROM32_INSTR_PT(589) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(601)
     OR ROM32_INSTR_PT(619) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(668) OR ROM32_INSTR_PT(674)
     OR ROM32_INSTR_PT(688) OR ROM32_INSTR_PT(694)
     OR ROM32_INSTR_PT(699) OR ROM32_INSTR_PT(702)
     OR ROM32_INSTR_PT(709) OR ROM32_INSTR_PT(714)
     OR ROM32_INSTR_PT(733) OR ROM32_INSTR_PT(778)
     OR ROM32_INSTR_PT(784) OR ROM32_INSTR_PT(812)
     OR ROM32_INSTR_PT(818) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(821) OR ROM32_INSTR_PT(824)
     OR ROM32_INSTR_PT(840) OR ROM32_INSTR_PT(843)
     OR ROM32_INSTR_PT(844) OR ROM32_INSTR_PT(847)
     OR ROM32_INSTR_PT(853) OR ROM32_INSTR_PT(878)
    );
MQQ1888:UCODE_END_EARLY <= 
    (ROM32_INSTR_PT(372) OR ROM32_INSTR_PT(389)
     OR ROM32_INSTR_PT(650) OR ROM32_INSTR_PT(673)
     OR ROM32_INSTR_PT(681) OR ROM32_INSTR_PT(687)
     OR ROM32_INSTR_PT(725) OR ROM32_INSTR_PT(734)
     OR ROM32_INSTR_PT(750) OR ROM32_INSTR_PT(754)
     OR ROM32_INSTR_PT(781) OR ROM32_INSTR_PT(782)
     OR ROM32_INSTR_PT(794) OR ROM32_INSTR_PT(796)
     OR ROM32_INSTR_PT(797) OR ROM32_INSTR_PT(802)
     OR ROM32_INSTR_PT(808) OR ROM32_INSTR_PT(813)
     OR ROM32_INSTR_PT(820) OR ROM32_INSTR_PT(827)
     OR ROM32_INSTR_PT(873));
MQQ1889:LOOP_BEGIN <= 
    (ROM32_INSTR_PT(24) OR ROM32_INSTR_PT(55)
     OR ROM32_INSTR_PT(105) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(147) OR ROM32_INSTR_PT(211)
     OR ROM32_INSTR_PT(228) OR ROM32_INSTR_PT(230)
     OR ROM32_INSTR_PT(239) OR ROM32_INSTR_PT(245)
     OR ROM32_INSTR_PT(253) OR ROM32_INSTR_PT(304)
     OR ROM32_INSTR_PT(308) OR ROM32_INSTR_PT(314)
     OR ROM32_INSTR_PT(321) OR ROM32_INSTR_PT(345)
     OR ROM32_INSTR_PT(366) OR ROM32_INSTR_PT(374)
     OR ROM32_INSTR_PT(407) OR ROM32_INSTR_PT(408)
     OR ROM32_INSTR_PT(432) OR ROM32_INSTR_PT(448)
     OR ROM32_INSTR_PT(460) OR ROM32_INSTR_PT(483)
     OR ROM32_INSTR_PT(490) OR ROM32_INSTR_PT(495)
     OR ROM32_INSTR_PT(544) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(571) OR ROM32_INSTR_PT(586)
     OR ROM32_INSTR_PT(604));
MQQ1890:LOOP_END <= 
    (ROM32_INSTR_PT(149) OR ROM32_INSTR_PT(156)
     OR ROM32_INSTR_PT(372) OR ROM32_INSTR_PT(466)
     OR ROM32_INSTR_PT(492) OR ROM32_INSTR_PT(500)
     OR ROM32_INSTR_PT(564) OR ROM32_INSTR_PT(637)
     OR ROM32_INSTR_PT(648) OR ROM32_INSTR_PT(655)
     OR ROM32_INSTR_PT(679) OR ROM32_INSTR_PT(696)
     OR ROM32_INSTR_PT(743) OR ROM32_INSTR_PT(769)
     OR ROM32_INSTR_PT(773) OR ROM32_INSTR_PT(783)
     OR ROM32_INSTR_PT(793) OR ROM32_INSTR_PT(802)
     OR ROM32_INSTR_PT(809) OR ROM32_INSTR_PT(810)
     OR ROM32_INSTR_PT(848) OR ROM32_INSTR_PT(861)
     OR ROM32_INSTR_PT(874));
MQQ1891:COUNT_SRC(0) <= 
    (ROM32_INSTR_PT(75) OR ROM32_INSTR_PT(744)
     OR ROM32_INSTR_PT(761) OR ROM32_INSTR_PT(875)
     OR ROM32_INSTR_PT(879) OR ROM32_INSTR_PT(880)
     OR ROM32_INSTR_PT(883) OR ROM32_INSTR_PT(890)
     OR ROM32_INSTR_PT(891) OR ROM32_INSTR_PT(892)
    );
MQQ1892:COUNT_SRC(1) <= 
    (ROM32_INSTR_PT(838) OR ROM32_INSTR_PT(875)
     OR ROM32_INSTR_PT(880) OR ROM32_INSTR_PT(882)
     OR ROM32_INSTR_PT(886) OR ROM32_INSTR_PT(891)
     OR ROM32_INSTR_PT(892));
MQQ1893:COUNT_SRC(2) <= 
    (ROM32_INSTR_PT(695) OR ROM32_INSTR_PT(744)
     OR ROM32_INSTR_PT(761) OR ROM32_INSTR_PT(828)
     OR ROM32_INSTR_PT(838) OR ROM32_INSTR_PT(890)
     OR ROM32_INSTR_PT(891) OR ROM32_INSTR_PT(892)
    );
MQQ1894:EXTRT <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(19)
     OR ROM32_INSTR_PT(21) OR ROM32_INSTR_PT(25)
     OR ROM32_INSTR_PT(40) OR ROM32_INSTR_PT(44)
     OR ROM32_INSTR_PT(47) OR ROM32_INSTR_PT(69)
     OR ROM32_INSTR_PT(72) OR ROM32_INSTR_PT(82)
     OR ROM32_INSTR_PT(91) OR ROM32_INSTR_PT(94)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(108)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(121)
     OR ROM32_INSTR_PT(131) OR ROM32_INSTR_PT(133)
     OR ROM32_INSTR_PT(136) OR ROM32_INSTR_PT(139)
     OR ROM32_INSTR_PT(151) OR ROM32_INSTR_PT(152)
     OR ROM32_INSTR_PT(161) OR ROM32_INSTR_PT(164)
     OR ROM32_INSTR_PT(168) OR ROM32_INSTR_PT(188)
     OR ROM32_INSTR_PT(190) OR ROM32_INSTR_PT(197)
     OR ROM32_INSTR_PT(221) OR ROM32_INSTR_PT(234)
     OR ROM32_INSTR_PT(236) OR ROM32_INSTR_PT(247)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(262)
     OR ROM32_INSTR_PT(265) OR ROM32_INSTR_PT(266)
     OR ROM32_INSTR_PT(277) OR ROM32_INSTR_PT(281)
     OR ROM32_INSTR_PT(284) OR ROM32_INSTR_PT(296)
     OR ROM32_INSTR_PT(300) OR ROM32_INSTR_PT(315)
     OR ROM32_INSTR_PT(316) OR ROM32_INSTR_PT(317)
     OR ROM32_INSTR_PT(327) OR ROM32_INSTR_PT(328)
     OR ROM32_INSTR_PT(333) OR ROM32_INSTR_PT(336)
     OR ROM32_INSTR_PT(349) OR ROM32_INSTR_PT(353)
     OR ROM32_INSTR_PT(354) OR ROM32_INSTR_PT(380)
     OR ROM32_INSTR_PT(381) OR ROM32_INSTR_PT(397)
     OR ROM32_INSTR_PT(410) OR ROM32_INSTR_PT(415)
     OR ROM32_INSTR_PT(420) OR ROM32_INSTR_PT(437)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(457)
     OR ROM32_INSTR_PT(461) OR ROM32_INSTR_PT(483)
     OR ROM32_INSTR_PT(493) OR ROM32_INSTR_PT(525)
     OR ROM32_INSTR_PT(529) OR ROM32_INSTR_PT(533)
     OR ROM32_INSTR_PT(536) OR ROM32_INSTR_PT(587)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(592)
     OR ROM32_INSTR_PT(594) OR ROM32_INSTR_PT(623)
     OR ROM32_INSTR_PT(627) OR ROM32_INSTR_PT(636)
     OR ROM32_INSTR_PT(645) OR ROM32_INSTR_PT(656)
     OR ROM32_INSTR_PT(665) OR ROM32_INSTR_PT(667)
     OR ROM32_INSTR_PT(669) OR ROM32_INSTR_PT(671)
     OR ROM32_INSTR_PT(686) OR ROM32_INSTR_PT(701)
     OR ROM32_INSTR_PT(707) OR ROM32_INSTR_PT(712)
     OR ROM32_INSTR_PT(721) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(723) OR ROM32_INSTR_PT(730)
     OR ROM32_INSTR_PT(735) OR ROM32_INSTR_PT(739)
     OR ROM32_INSTR_PT(742) OR ROM32_INSTR_PT(746)
     OR ROM32_INSTR_PT(756) OR ROM32_INSTR_PT(757)
     OR ROM32_INSTR_PT(758) OR ROM32_INSTR_PT(760)
     OR ROM32_INSTR_PT(764) OR ROM32_INSTR_PT(765)
     OR ROM32_INSTR_PT(766) OR ROM32_INSTR_PT(767)
     OR ROM32_INSTR_PT(768) OR ROM32_INSTR_PT(771)
     OR ROM32_INSTR_PT(772) OR ROM32_INSTR_PT(775)
     OR ROM32_INSTR_PT(776) OR ROM32_INSTR_PT(777)
     OR ROM32_INSTR_PT(788) OR ROM32_INSTR_PT(789)
     OR ROM32_INSTR_PT(791) OR ROM32_INSTR_PT(792)
     OR ROM32_INSTR_PT(798) OR ROM32_INSTR_PT(804)
     OR ROM32_INSTR_PT(806) OR ROM32_INSTR_PT(811)
     OR ROM32_INSTR_PT(816) OR ROM32_INSTR_PT(826)
     OR ROM32_INSTR_PT(833) OR ROM32_INSTR_PT(834)
     OR ROM32_INSTR_PT(835) OR ROM32_INSTR_PT(837)
     OR ROM32_INSTR_PT(841) OR ROM32_INSTR_PT(849)
     OR ROM32_INSTR_PT(856) OR ROM32_INSTR_PT(858)
     OR ROM32_INSTR_PT(859) OR ROM32_INSTR_PT(860)
     OR ROM32_INSTR_PT(862) OR ROM32_INSTR_PT(863)
     OR ROM32_INSTR_PT(864) OR ROM32_INSTR_PT(865)
     OR ROM32_INSTR_PT(866) OR ROM32_INSTR_PT(867)
     OR ROM32_INSTR_PT(870) OR ROM32_INSTR_PT(876)
     OR ROM32_INSTR_PT(884) OR ROM32_INSTR_PT(885)
    );
MQQ1895:EXTS1 <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(19)
     OR ROM32_INSTR_PT(21) OR ROM32_INSTR_PT(28)
     OR ROM32_INSTR_PT(36) OR ROM32_INSTR_PT(47)
     OR ROM32_INSTR_PT(58) OR ROM32_INSTR_PT(82)
     OR ROM32_INSTR_PT(91) OR ROM32_INSTR_PT(100)
     OR ROM32_INSTR_PT(107) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(136) OR ROM32_INSTR_PT(137)
     OR ROM32_INSTR_PT(157) OR ROM32_INSTR_PT(167)
     OR ROM32_INSTR_PT(193) OR ROM32_INSTR_PT(197)
     OR ROM32_INSTR_PT(212) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(231) OR ROM32_INSTR_PT(236)
     OR ROM32_INSTR_PT(263) OR ROM32_INSTR_PT(277)
     OR ROM32_INSTR_PT(286) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(296) OR ROM32_INSTR_PT(298)
     OR ROM32_INSTR_PT(315) OR ROM32_INSTR_PT(316)
     OR ROM32_INSTR_PT(317) OR ROM32_INSTR_PT(324)
     OR ROM32_INSTR_PT(327) OR ROM32_INSTR_PT(328)
     OR ROM32_INSTR_PT(330) OR ROM32_INSTR_PT(336)
     OR ROM32_INSTR_PT(346) OR ROM32_INSTR_PT(369)
     OR ROM32_INSTR_PT(380) OR ROM32_INSTR_PT(397)
     OR ROM32_INSTR_PT(410) OR ROM32_INSTR_PT(414)
     OR ROM32_INSTR_PT(438) OR ROM32_INSTR_PT(447)
     OR ROM32_INSTR_PT(457) OR ROM32_INSTR_PT(462)
     OR ROM32_INSTR_PT(470) OR ROM32_INSTR_PT(488)
     OR ROM32_INSTR_PT(493) OR ROM32_INSTR_PT(495)
     OR ROM32_INSTR_PT(499) OR ROM32_INSTR_PT(526)
     OR ROM32_INSTR_PT(542) OR ROM32_INSTR_PT(589)
     OR ROM32_INSTR_PT(594) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(623) OR ROM32_INSTR_PT(627)
     OR ROM32_INSTR_PT(636) OR ROM32_INSTR_PT(645)
     OR ROM32_INSTR_PT(651) OR ROM32_INSTR_PT(656)
     OR ROM32_INSTR_PT(667) OR ROM32_INSTR_PT(669)
     OR ROM32_INSTR_PT(670) OR ROM32_INSTR_PT(675)
     OR ROM32_INSTR_PT(686) OR ROM32_INSTR_PT(691)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(701)
     OR ROM32_INSTR_PT(706) OR ROM32_INSTR_PT(707)
     OR ROM32_INSTR_PT(710) OR ROM32_INSTR_PT(716)
     OR ROM32_INSTR_PT(721) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(730) OR ROM32_INSTR_PT(733)
     OR ROM32_INSTR_PT(739) OR ROM32_INSTR_PT(741)
     OR ROM32_INSTR_PT(742) OR ROM32_INSTR_PT(746)
     OR ROM32_INSTR_PT(756) OR ROM32_INSTR_PT(757)
     OR ROM32_INSTR_PT(758) OR ROM32_INSTR_PT(760)
     OR ROM32_INSTR_PT(764) OR ROM32_INSTR_PT(765)
     OR ROM32_INSTR_PT(767) OR ROM32_INSTR_PT(768)
     OR ROM32_INSTR_PT(771) OR ROM32_INSTR_PT(775)
     OR ROM32_INSTR_PT(776) OR ROM32_INSTR_PT(777)
     OR ROM32_INSTR_PT(779) OR ROM32_INSTR_PT(788)
     OR ROM32_INSTR_PT(789) OR ROM32_INSTR_PT(791)
     OR ROM32_INSTR_PT(798) OR ROM32_INSTR_PT(801)
     OR ROM32_INSTR_PT(804) OR ROM32_INSTR_PT(806)
     OR ROM32_INSTR_PT(811) OR ROM32_INSTR_PT(812)
     OR ROM32_INSTR_PT(816) OR ROM32_INSTR_PT(824)
     OR ROM32_INSTR_PT(826) OR ROM32_INSTR_PT(830)
     OR ROM32_INSTR_PT(832) OR ROM32_INSTR_PT(833)
     OR ROM32_INSTR_PT(835) OR ROM32_INSTR_PT(837)
     OR ROM32_INSTR_PT(841) OR ROM32_INSTR_PT(842)
     OR ROM32_INSTR_PT(843) OR ROM32_INSTR_PT(846)
     OR ROM32_INSTR_PT(847) OR ROM32_INSTR_PT(849)
     OR ROM32_INSTR_PT(850) OR ROM32_INSTR_PT(852)
     OR ROM32_INSTR_PT(858) OR ROM32_INSTR_PT(859)
     OR ROM32_INSTR_PT(863) OR ROM32_INSTR_PT(865)
     OR ROM32_INSTR_PT(867) OR ROM32_INSTR_PT(868)
     OR ROM32_INSTR_PT(877) OR ROM32_INSTR_PT(878)
     OR ROM32_INSTR_PT(888));
MQQ1896:EXTS2 <= 
    (ROM32_INSTR_PT(21) OR ROM32_INSTR_PT(25)
     OR ROM32_INSTR_PT(36) OR ROM32_INSTR_PT(44)
     OR ROM32_INSTR_PT(47) OR ROM32_INSTR_PT(91)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(136)
     OR ROM32_INSTR_PT(137) OR ROM32_INSTR_PT(139)
     OR ROM32_INSTR_PT(152) OR ROM32_INSTR_PT(167)
     OR ROM32_INSTR_PT(178) OR ROM32_INSTR_PT(188)
     OR ROM32_INSTR_PT(191) OR ROM32_INSTR_PT(212)
     OR ROM32_INSTR_PT(217) OR ROM32_INSTR_PT(236)
     OR ROM32_INSTR_PT(295) OR ROM32_INSTR_PT(317)
     OR ROM32_INSTR_PT(327) OR ROM32_INSTR_PT(328)
     OR ROM32_INSTR_PT(330) OR ROM32_INSTR_PT(333)
     OR ROM32_INSTR_PT(336) OR ROM32_INSTR_PT(341)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(346)
     OR ROM32_INSTR_PT(354) OR ROM32_INSTR_PT(356)
     OR ROM32_INSTR_PT(369) OR ROM32_INSTR_PT(375)
     OR ROM32_INSTR_PT(381) OR ROM32_INSTR_PT(393)
     OR ROM32_INSTR_PT(410) OR ROM32_INSTR_PT(415)
     OR ROM32_INSTR_PT(429) OR ROM32_INSTR_PT(437)
     OR ROM32_INSTR_PT(438) OR ROM32_INSTR_PT(447)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(457)
     OR ROM32_INSTR_PT(470) OR ROM32_INSTR_PT(493)
     OR ROM32_INSTR_PT(518) OR ROM32_INSTR_PT(526)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(579)
     OR ROM32_INSTR_PT(587) OR ROM32_INSTR_PT(594)
     OR ROM32_INSTR_PT(599) OR ROM32_INSTR_PT(624)
     OR ROM32_INSTR_PT(627) OR ROM32_INSTR_PT(628)
     OR ROM32_INSTR_PT(651) OR ROM32_INSTR_PT(656)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(706)
     OR ROM32_INSTR_PT(710) OR ROM32_INSTR_PT(714)
     OR ROM32_INSTR_PT(721) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(723) OR ROM32_INSTR_PT(730)
     OR ROM32_INSTR_PT(735) OR ROM32_INSTR_PT(737)
     OR ROM32_INSTR_PT(739) OR ROM32_INSTR_PT(742)
     OR ROM32_INSTR_PT(746) OR ROM32_INSTR_PT(749)
     OR ROM32_INSTR_PT(756) OR ROM32_INSTR_PT(760)
     OR ROM32_INSTR_PT(764) OR ROM32_INSTR_PT(767)
     OR ROM32_INSTR_PT(770) OR ROM32_INSTR_PT(779)
     OR ROM32_INSTR_PT(789) OR ROM32_INSTR_PT(791)
     OR ROM32_INSTR_PT(812) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(822) OR ROM32_INSTR_PT(824)
     OR ROM32_INSTR_PT(835) OR ROM32_INSTR_PT(841)
     OR ROM32_INSTR_PT(842) OR ROM32_INSTR_PT(850)
     OR ROM32_INSTR_PT(853) OR ROM32_INSTR_PT(858)
     OR ROM32_INSTR_PT(863) OR ROM32_INSTR_PT(865)
     OR ROM32_INSTR_PT(867) OR ROM32_INSTR_PT(868)
     OR ROM32_INSTR_PT(876) OR ROM32_INSTR_PT(878)
     OR ROM32_INSTR_PT(885));
MQQ1897:EXTS3 <= 
    (ROM32_INSTR_PT(47) OR ROM32_INSTR_PT(58)
     OR ROM32_INSTR_PT(126) OR ROM32_INSTR_PT(133)
     OR ROM32_INSTR_PT(135) OR ROM32_INSTR_PT(168)
     OR ROM32_INSTR_PT(190) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(263) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(333)
     OR ROM32_INSTR_PT(346) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(397) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(467) OR ROM32_INSTR_PT(487)
     OR ROM32_INSTR_PT(526) OR ROM32_INSTR_PT(623)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(707)
     OR ROM32_INSTR_PT(710) OR ROM32_INSTR_PT(717)
     OR ROM32_INSTR_PT(730) OR ROM32_INSTR_PT(771)
     OR ROM32_INSTR_PT(792) OR ROM32_INSTR_PT(804)
     OR ROM32_INSTR_PT(826) OR ROM32_INSTR_PT(837)
     OR ROM32_INSTR_PT(866) OR ROM32_INSTR_PT(887)
    );
MQQ1898:SEL0_5 <= 
    (ROM32_INSTR_PT(651) OR ROM32_INSTR_PT(714)
    );
MQQ1899:SEL6_10(0) <= 
    (ROM32_INSTR_PT(40) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(83) OR ROM32_INSTR_PT(94)
     OR ROM32_INSTR_PT(108) OR ROM32_INSTR_PT(201)
     OR ROM32_INSTR_PT(212) OR ROM32_INSTR_PT(266)
     OR ROM32_INSTR_PT(384) OR ROM32_INSTR_PT(438)
     OR ROM32_INSTR_PT(440) OR ROM32_INSTR_PT(450)
     OR ROM32_INSTR_PT(512) OR ROM32_INSTR_PT(518)
     OR ROM32_INSTR_PT(528) OR ROM32_INSTR_PT(529)
     OR ROM32_INSTR_PT(536) OR ROM32_INSTR_PT(541)
     OR ROM32_INSTR_PT(548) OR ROM32_INSTR_PT(559)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(572)
     OR ROM32_INSTR_PT(580) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(601) OR ROM32_INSTR_PT(618)
     OR ROM32_INSTR_PT(661) OR ROM32_INSTR_PT(693)
     OR ROM32_INSTR_PT(702) OR ROM32_INSTR_PT(784)
     OR ROM32_INSTR_PT(818) OR ROM32_INSTR_PT(853)
    );
MQQ1900:SEL6_10(1) <= 
    (ROM32_INSTR_PT(1) OR ROM32_INSTR_PT(2)
     OR ROM32_INSTR_PT(40) OR ROM32_INSTR_PT(54)
     OR ROM32_INSTR_PT(71) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(80) OR ROM32_INSTR_PT(83)
     OR ROM32_INSTR_PT(94) OR ROM32_INSTR_PT(108)
     OR ROM32_INSTR_PT(121) OR ROM32_INSTR_PT(178)
     OR ROM32_INSTR_PT(182) OR ROM32_INSTR_PT(262)
     OR ROM32_INSTR_PT(266) OR ROM32_INSTR_PT(284)
     OR ROM32_INSTR_PT(334) OR ROM32_INSTR_PT(344)
     OR ROM32_INSTR_PT(346) OR ROM32_INSTR_PT(347)
     OR ROM32_INSTR_PT(351) OR ROM32_INSTR_PT(356)
     OR ROM32_INSTR_PT(375) OR ROM32_INSTR_PT(403)
     OR ROM32_INSTR_PT(427) OR ROM32_INSTR_PT(432)
     OR ROM32_INSTR_PT(455) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(483) OR ROM32_INSTR_PT(485)
     OR ROM32_INSTR_PT(529) OR ROM32_INSTR_PT(530)
     OR ROM32_INSTR_PT(536) OR ROM32_INSTR_PT(539)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(592)
     OR ROM32_INSTR_PT(651) OR ROM32_INSTR_PT(658)
     OR ROM32_INSTR_PT(691) OR ROM32_INSTR_PT(692)
     OR ROM32_INSTR_PT(703) OR ROM32_INSTR_PT(710)
     OR ROM32_INSTR_PT(714) OR ROM32_INSTR_PT(716)
     OR ROM32_INSTR_PT(723) OR ROM32_INSTR_PT(724)
     OR ROM32_INSTR_PT(732) OR ROM32_INSTR_PT(856)
     OR ROM32_INSTR_PT(862) OR ROM32_INSTR_PT(870)
    );
MQQ1901:SEL11_15(0) <= 
    (ROM32_INSTR_PT(36) OR ROM32_INSTR_PT(133)
     OR ROM32_INSTR_PT(193) OR ROM32_INSTR_PT(231)
     OR ROM32_INSTR_PT(246) OR ROM32_INSTR_PT(286)
     OR ROM32_INSTR_PT(369) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(444)
     OR ROM32_INSTR_PT(462) OR ROM32_INSTR_PT(589)
     OR ROM32_INSTR_PT(663) OR ROM32_INSTR_PT(733)
     OR ROM32_INSTR_PT(792) OR ROM32_INSTR_PT(825)
    );
MQQ1902:SEL11_15(1) <= 
    (ROM32_INSTR_PT(22) OR ROM32_INSTR_PT(25)
     OR ROM32_INSTR_PT(36) OR ROM32_INSTR_PT(44)
     OR ROM32_INSTR_PT(48) OR ROM32_INSTR_PT(61)
     OR ROM32_INSTR_PT(64) OR ROM32_INSTR_PT(65)
     OR ROM32_INSTR_PT(69) OR ROM32_INSTR_PT(86)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(106)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(129)
     OR ROM32_INSTR_PT(131) OR ROM32_INSTR_PT(139)
     OR ROM32_INSTR_PT(140) OR ROM32_INSTR_PT(151)
     OR ROM32_INSTR_PT(160) OR ROM32_INSTR_PT(164)
     OR ROM32_INSTR_PT(188) OR ROM32_INSTR_PT(190)
     OR ROM32_INSTR_PT(193) OR ROM32_INSTR_PT(201)
     OR ROM32_INSTR_PT(221) OR ROM32_INSTR_PT(231)
     OR ROM32_INSTR_PT(234) OR ROM32_INSTR_PT(247)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(265)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(286)
     OR ROM32_INSTR_PT(300) OR ROM32_INSTR_PT(351)
     OR ROM32_INSTR_PT(354) OR ROM32_INSTR_PT(369)
     OR ROM32_INSTR_PT(384) OR ROM32_INSTR_PT(393)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(420)
     OR ROM32_INSTR_PT(429) OR ROM32_INSTR_PT(434)
     OR ROM32_INSTR_PT(437) OR ROM32_INSTR_PT(440)
     OR ROM32_INSTR_PT(450) OR ROM32_INSTR_PT(451)
     OR ROM32_INSTR_PT(462) OR ROM32_INSTR_PT(518)
     OR ROM32_INSTR_PT(523) OR ROM32_INSTR_PT(528)
     OR ROM32_INSTR_PT(545) OR ROM32_INSTR_PT(548)
     OR ROM32_INSTR_PT(559) OR ROM32_INSTR_PT(572)
     OR ROM32_INSTR_PT(587) OR ROM32_INSTR_PT(589)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(601)
     OR ROM32_INSTR_PT(618) OR ROM32_INSTR_PT(624)
     OR ROM32_INSTR_PT(631) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(665) OR ROM32_INSTR_PT(693)
     OR ROM32_INSTR_PT(702) OR ROM32_INSTR_PT(713)
     OR ROM32_INSTR_PT(714) OR ROM32_INSTR_PT(727)
     OR ROM32_INSTR_PT(780) OR ROM32_INSTR_PT(784)
     OR ROM32_INSTR_PT(801) OR ROM32_INSTR_PT(812)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(824)
     OR ROM32_INSTR_PT(839) OR ROM32_INSTR_PT(843)
     OR ROM32_INSTR_PT(847) OR ROM32_INSTR_PT(878)
    );
MQQ1903:SEL16_20(0) <= 
    (ROM32_INSTR_PT(5) OR ROM32_INSTR_PT(133)
     OR ROM32_INSTR_PT(194) OR ROM32_INSTR_PT(254)
     OR ROM32_INSTR_PT(256) OR ROM32_INSTR_PT(353)
     OR ROM32_INSTR_PT(444) OR ROM32_INSTR_PT(533)
     OR ROM32_INSTR_PT(792) OR ROM32_INSTR_PT(825)
    );
MQQ1904:SEL16_20(1) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(11)
     OR ROM32_INSTR_PT(15) OR ROM32_INSTR_PT(28)
     OR ROM32_INSTR_PT(40) OR ROM32_INSTR_PT(46)
     OR ROM32_INSTR_PT(48) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(76) OR ROM32_INSTR_PT(83)
     OR ROM32_INSTR_PT(88) OR ROM32_INSTR_PT(94)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(108)
     OR ROM32_INSTR_PT(126) OR ROM32_INSTR_PT(131)
     OR ROM32_INSTR_PT(133) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(140) OR ROM32_INSTR_PT(161)
     OR ROM32_INSTR_PT(164) OR ROM32_INSTR_PT(201)
     OR ROM32_INSTR_PT(204) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(248) OR ROM32_INSTR_PT(265)
     OR ROM32_INSTR_PT(266) OR ROM32_INSTR_PT(277)
     OR ROM32_INSTR_PT(293) OR ROM32_INSTR_PT(298)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(320)
     OR ROM32_INSTR_PT(334) OR ROM32_INSTR_PT(351)
     OR ROM32_INSTR_PT(353) OR ROM32_INSTR_PT(359)
     OR ROM32_INSTR_PT(384) OR ROM32_INSTR_PT(397)
     OR ROM32_INSTR_PT(409) OR ROM32_INSTR_PT(420)
     OR ROM32_INSTR_PT(443) OR ROM32_INSTR_PT(444)
     OR ROM32_INSTR_PT(450) OR ROM32_INSTR_PT(467)
     OR ROM32_INSTR_PT(487) OR ROM32_INSTR_PT(495)
     OR ROM32_INSTR_PT(510) OR ROM32_INSTR_PT(523)
     OR ROM32_INSTR_PT(528) OR ROM32_INSTR_PT(529)
     OR ROM32_INSTR_PT(540) OR ROM32_INSTR_PT(548)
     OR ROM32_INSTR_PT(559) OR ROM32_INSTR_PT(560)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(571)
     OR ROM32_INSTR_PT(572) OR ROM32_INSTR_PT(600)
     OR ROM32_INSTR_PT(601) OR ROM32_INSTR_PT(609)
     OR ROM32_INSTR_PT(618) OR ROM32_INSTR_PT(631)
     OR ROM32_INSTR_PT(649) OR ROM32_INSTR_PT(661)
     OR ROM32_INSTR_PT(693) OR ROM32_INSTR_PT(702)
     OR ROM32_INSTR_PT(713) OR ROM32_INSTR_PT(766)
     OR ROM32_INSTR_PT(784) OR ROM32_INSTR_PT(792)
     OR ROM32_INSTR_PT(825) OR ROM32_INSTR_PT(836)
    );
MQQ1905:SEL21_25(0) <= 
    (ROM32_INSTR_PT(197));
MQQ1906:SEL21_25(1) <= 
    (ROM32_INSTR_PT(15) OR ROM32_INSTR_PT(28)
     OR ROM32_INSTR_PT(46) OR ROM32_INSTR_PT(48)
     OR ROM32_INSTR_PT(65) OR ROM32_INSTR_PT(76)
     OR ROM32_INSTR_PT(88) OR ROM32_INSTR_PT(140)
     OR ROM32_INSTR_PT(201) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(265) OR ROM32_INSTR_PT(320)
     OR ROM32_INSTR_PT(351) OR ROM32_INSTR_PT(359)
     OR ROM32_INSTR_PT(384) OR ROM32_INSTR_PT(420)
     OR ROM32_INSTR_PT(450) OR ROM32_INSTR_PT(467)
     OR ROM32_INSTR_PT(512) OR ROM32_INSTR_PT(528)
     OR ROM32_INSTR_PT(540) OR ROM32_INSTR_PT(548)
     OR ROM32_INSTR_PT(559) OR ROM32_INSTR_PT(571)
     OR ROM32_INSTR_PT(572) OR ROM32_INSTR_PT(631)
     OR ROM32_INSTR_PT(651) OR ROM32_INSTR_PT(702)
     OR ROM32_INSTR_PT(714) OR ROM32_INSTR_PT(727)
     OR ROM32_INSTR_PT(784));
MQQ1907:SEL26_30 <= 
    (ROM32_INSTR_PT(15) OR ROM32_INSTR_PT(28)
     OR ROM32_INSTR_PT(46) OR ROM32_INSTR_PT(48)
     OR ROM32_INSTR_PT(65) OR ROM32_INSTR_PT(76)
     OR ROM32_INSTR_PT(88) OR ROM32_INSTR_PT(140)
     OR ROM32_INSTR_PT(201) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(265) OR ROM32_INSTR_PT(320)
     OR ROM32_INSTR_PT(351) OR ROM32_INSTR_PT(359)
     OR ROM32_INSTR_PT(384) OR ROM32_INSTR_PT(420)
     OR ROM32_INSTR_PT(450) OR ROM32_INSTR_PT(467)
     OR ROM32_INSTR_PT(512) OR ROM32_INSTR_PT(528)
     OR ROM32_INSTR_PT(540) OR ROM32_INSTR_PT(548)
     OR ROM32_INSTR_PT(559) OR ROM32_INSTR_PT(571)
     OR ROM32_INSTR_PT(572) OR ROM32_INSTR_PT(631)
     OR ROM32_INSTR_PT(651) OR ROM32_INSTR_PT(702)
     OR ROM32_INSTR_PT(714) OR ROM32_INSTR_PT(727)
     OR ROM32_INSTR_PT(784));
MQQ1908:SEL31 <= 
    (ROM32_INSTR_PT(15) OR ROM32_INSTR_PT(28)
     OR ROM32_INSTR_PT(61) OR ROM32_INSTR_PT(65)
     OR ROM32_INSTR_PT(76) OR ROM32_INSTR_PT(88)
     OR ROM32_INSTR_PT(140) OR ROM32_INSTR_PT(201)
     OR ROM32_INSTR_PT(265) OR ROM32_INSTR_PT(320)
     OR ROM32_INSTR_PT(346) OR ROM32_INSTR_PT(351)
     OR ROM32_INSTR_PT(356) OR ROM32_INSTR_PT(359)
     OR ROM32_INSTR_PT(384) OR ROM32_INSTR_PT(420)
     OR ROM32_INSTR_PT(450) OR ROM32_INSTR_PT(467)
     OR ROM32_INSTR_PT(540) OR ROM32_INSTR_PT(541)
     OR ROM32_INSTR_PT(559) OR ROM32_INSTR_PT(560)
     OR ROM32_INSTR_PT(572) OR ROM32_INSTR_PT(631)
     OR ROM32_INSTR_PT(651) OR ROM32_INSTR_PT(692)
     OR ROM32_INSTR_PT(702) OR ROM32_INSTR_PT(710)
     OR ROM32_INSTR_PT(714) OR ROM32_INSTR_PT(784)
     OR ROM32_INSTR_PT(818));
MQQ1909:CR_BF2FXM <= 
    (ROM32_INSTR_PT(713));
MQQ1910:SKIP_COND <= 
    (ROM32_INSTR_PT(21) OR ROM32_INSTR_PT(32)
     OR ROM32_INSTR_PT(82) OR ROM32_INSTR_PT(89)
     OR ROM32_INSTR_PT(91) OR ROM32_INSTR_PT(127)
     OR ROM32_INSTR_PT(217) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(327) OR ROM32_INSTR_PT(328)
     OR ROM32_INSTR_PT(341) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(485) OR ROM32_INSTR_PT(662)
     OR ROM32_INSTR_PT(667) OR ROM32_INSTR_PT(676)
     OR ROM32_INSTR_PT(682) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(736) OR ROM32_INSTR_PT(737)
     OR ROM32_INSTR_PT(738) OR ROM32_INSTR_PT(739)
     OR ROM32_INSTR_PT(740) OR ROM32_INSTR_PT(742)
     OR ROM32_INSTR_PT(747) OR ROM32_INSTR_PT(748)
     OR ROM32_INSTR_PT(749) OR ROM32_INSTR_PT(758)
     OR ROM32_INSTR_PT(770) OR ROM32_INSTR_PT(775)
     OR ROM32_INSTR_PT(776) OR ROM32_INSTR_PT(777)
     OR ROM32_INSTR_PT(786) OR ROM32_INSTR_PT(788)
     OR ROM32_INSTR_PT(789) OR ROM32_INSTR_PT(800)
     OR ROM32_INSTR_PT(811) OR ROM32_INSTR_PT(814)
     OR ROM32_INSTR_PT(815) OR ROM32_INSTR_PT(816)
     OR ROM32_INSTR_PT(822) OR ROM32_INSTR_PT(842)
     OR ROM32_INSTR_PT(858) OR ROM32_INSTR_PT(865)
    );
MQQ1911:SKIP_ZERO <= 
    (ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(349)
     OR ROM32_INSTR_PT(432) OR ROM32_INSTR_PT(457)
     OR ROM32_INSTR_PT(483) OR ROM32_INSTR_PT(671)
     OR ROM32_INSTR_PT(712));
MQQ1912:LOOP_ADDR(0) <= 
    (ROM32_INSTR_PT(19) OR ROM32_INSTR_PT(36)
     OR ROM32_INSTR_PT(58) OR ROM32_INSTR_PT(315)
     OR ROM32_INSTR_PT(316) OR ROM32_INSTR_PT(349)
     OR ROM32_INSTR_PT(369) OR ROM32_INSTR_PT(457)
     OR ROM32_INSTR_PT(623) OR ROM32_INSTR_PT(627)
     OR ROM32_INSTR_PT(656) OR ROM32_INSTR_PT(671)
     OR ROM32_INSTR_PT(712) OR ROM32_INSTR_PT(721)
     OR ROM32_INSTR_PT(730) OR ROM32_INSTR_PT(742)
     OR ROM32_INSTR_PT(760) OR ROM32_INSTR_PT(771)
     OR ROM32_INSTR_PT(777) OR ROM32_INSTR_PT(798)
     OR ROM32_INSTR_PT(837) OR ROM32_INSTR_PT(863)
     OR ROM32_INSTR_PT(865));
MQQ1913:LOOP_ADDR(1) <= 
    (ROM32_INSTR_PT(315) OR ROM32_INSTR_PT(525)
     OR ROM32_INSTR_PT(623) OR ROM32_INSTR_PT(627)
     OR ROM32_INSTR_PT(656) OR ROM32_INSTR_PT(712)
     OR ROM32_INSTR_PT(721) OR ROM32_INSTR_PT(730)
     OR ROM32_INSTR_PT(742) OR ROM32_INSTR_PT(777)
     OR ROM32_INSTR_PT(837) OR ROM32_INSTR_PT(858)
     OR ROM32_INSTR_PT(865));
MQQ1914:LOOP_ADDR(2) <= 
    (ROM32_INSTR_PT(58) OR ROM32_INSTR_PT(457)
     OR ROM32_INSTR_PT(717) OR ROM32_INSTR_PT(740)
     OR ROM32_INSTR_PT(747) OR ROM32_INSTR_PT(887)
    );
MQQ1915:LOOP_ADDR(3) <= 
    (ROM32_INSTR_PT(19) OR ROM32_INSTR_PT(58)
     OR ROM32_INSTR_PT(136) OR ROM32_INSTR_PT(316)
     OR ROM32_INSTR_PT(414) OR ROM32_INSTR_PT(457)
     OR ROM32_INSTR_PT(623) OR ROM32_INSTR_PT(706)
     OR ROM32_INSTR_PT(722) OR ROM32_INSTR_PT(730)
     OR ROM32_INSTR_PT(756) OR ROM32_INSTR_PT(760)
     OR ROM32_INSTR_PT(771) OR ROM32_INSTR_PT(798)
     OR ROM32_INSTR_PT(837) OR ROM32_INSTR_PT(864)
     OR ROM32_INSTR_PT(865));
MQQ1916:LOOP_ADDR(4) <= 
    (ROM32_INSTR_PT(19) OR ROM32_INSTR_PT(36)
     OR ROM32_INSTR_PT(58) OR ROM32_INSTR_PT(136)
     OR ROM32_INSTR_PT(315) OR ROM32_INSTR_PT(349)
     OR ROM32_INSTR_PT(369) OR ROM32_INSTR_PT(410)
     OR ROM32_INSTR_PT(457) OR ROM32_INSTR_PT(470)
     OR ROM32_INSTR_PT(717) OR ROM32_INSTR_PT(740)
     OR ROM32_INSTR_PT(742) OR ROM32_INSTR_PT(747)
     OR ROM32_INSTR_PT(777) OR ROM32_INSTR_PT(837)
     OR ROM32_INSTR_PT(863) OR ROM32_INSTR_PT(865)
    );
MQQ1917:LOOP_ADDR(5) <= 
    (ROM32_INSTR_PT(36) OR ROM32_INSTR_PT(58)
     OR ROM32_INSTR_PT(315) OR ROM32_INSTR_PT(623)
     OR ROM32_INSTR_PT(656) OR ROM32_INSTR_PT(671)
     OR ROM32_INSTR_PT(721) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(735) OR ROM32_INSTR_PT(756)
     OR ROM32_INSTR_PT(764) OR ROM32_INSTR_PT(771)
     OR ROM32_INSTR_PT(798) OR ROM32_INSTR_PT(863)
    );
MQQ1918:LOOP_ADDR(6) <= 
    (ROM32_INSTR_PT(36) OR ROM32_INSTR_PT(136)
     OR ROM32_INSTR_PT(315) OR ROM32_INSTR_PT(316)
     OR ROM32_INSTR_PT(369) OR ROM32_INSTR_PT(380)
     OR ROM32_INSTR_PT(457) OR ROM32_INSTR_PT(470)
     OR ROM32_INSTR_PT(623) OR ROM32_INSTR_PT(671)
     OR ROM32_INSTR_PT(721) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(740) OR ROM32_INSTR_PT(742)
     OR ROM32_INSTR_PT(756) OR ROM32_INSTR_PT(760)
     OR ROM32_INSTR_PT(837) OR ROM32_INSTR_PT(858)
     OR ROM32_INSTR_PT(887));
MQQ1919:LOOP_ADDR(7) <= 
    (ROM32_INSTR_PT(19) OR ROM32_INSTR_PT(36)
     OR ROM32_INSTR_PT(58) OR ROM32_INSTR_PT(316)
     OR ROM32_INSTR_PT(349) OR ROM32_INSTR_PT(380)
     OR ROM32_INSTR_PT(410) OR ROM32_INSTR_PT(414)
     OR ROM32_INSTR_PT(623) OR ROM32_INSTR_PT(627)
     OR ROM32_INSTR_PT(721) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(730) OR ROM32_INSTR_PT(740)
     OR ROM32_INSTR_PT(742) OR ROM32_INSTR_PT(765)
     OR ROM32_INSTR_PT(771) OR ROM32_INSTR_PT(826)
     OR ROM32_INSTR_PT(865));
MQQ1920:LOOP_ADDR(8) <= 
    (ROM32_INSTR_PT(136) OR ROM32_INSTR_PT(410)
     OR ROM32_INSTR_PT(414) OR ROM32_INSTR_PT(457)
     OR ROM32_INSTR_PT(470) OR ROM32_INSTR_PT(488)
     OR ROM32_INSTR_PT(706) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(730) OR ROM32_INSTR_PT(740)
     OR ROM32_INSTR_PT(742) OR ROM32_INSTR_PT(747)
     OR ROM32_INSTR_PT(756) OR ROM32_INSTR_PT(863)
     OR ROM32_INSTR_PT(887));
MQQ1921:LOOP_ADDR(9) <= 
    (ROM32_INSTR_PT(19) OR ROM32_INSTR_PT(36)
     OR ROM32_INSTR_PT(58) OR ROM32_INSTR_PT(191)
     OR ROM32_INSTR_PT(316) OR ROM32_INSTR_PT(349)
     OR ROM32_INSTR_PT(369) OR ROM32_INSTR_PT(525)
     OR ROM32_INSTR_PT(623) OR ROM32_INSTR_PT(671)
     OR ROM32_INSTR_PT(717) OR ROM32_INSTR_PT(721)
     OR ROM32_INSTR_PT(760) OR ROM32_INSTR_PT(771)
     OR ROM32_INSTR_PT(777) OR ROM32_INSTR_PT(837)
     OR ROM32_INSTR_PT(887));
MQQ1922:LOOP_INIT(0) <= 
    (ROM32_INSTR_PT(168) OR ROM32_INSTR_PT(236)
     OR ROM32_INSTR_PT(315) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(397) OR ROM32_INSTR_PT(686)
     OR ROM32_INSTR_PT(717) OR ROM32_INSTR_PT(776)
     OR ROM32_INSTR_PT(788) OR ROM32_INSTR_PT(811)
     OR ROM32_INSTR_PT(816) OR ROM32_INSTR_PT(864)
    );
MQQ1923:LOOP_INIT(1) <= 
    (ROM32_INSTR_PT(893));
MQQ1924:LOOP_INIT(2) <= 
    (ROM32_INSTR_PT(168) OR ROM32_INSTR_PT(776)
     OR ROM32_INSTR_PT(811));
MQQ1925:EP <= 
    (ROM32_INSTR_PT(44) OR ROM32_INSTR_PT(61)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(277) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(354) OR ROM32_INSTR_PT(393)
     OR ROM32_INSTR_PT(397) OR ROM32_INSTR_PT(429)
     OR ROM32_INSTR_PT(437) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(523) OR ROM32_INSTR_PT(560)
    );

end generate;
rom_addr_d  <=  rom_addr;
rom_data  <=  template & ucode_end & ucode_end_early & loop_begin & loop_end & count_src & extRT & extS1 & extS2 & extS3 &
            sel0_5 & sel6_10 & sel11_15 & sel16_20 & sel21_25 & sel26_30 & sel31 & cr_bf2fxm & skip_cond & skip_zero & loop_addr & loop_init & ep;
-----------------------------------------------------------------------
-- Latches
-----------------------------------------------------------------------
rom_addr_latch: tri_rlmreg_p
  generic map (width => rom_addr_l2'length, init => 0, needs_sreset => 0, expand_type => expand_type)
  port map (vd      => vdd,
            gd      => gnd,
            nclk    => nclk,
            act     => rom_act,
            thold_b => pc_iu_func_sl_thold_0_b,
            sg      => pc_iu_sg_0,
            forcee => forcee,
            delay_lclkr => delay_lclkr,
            mpw1_b      => mpw1_b,
            mpw2_b      => mpw2_b,
            d_mode      => d_mode,
            scin    => siv(rom_addr_offset to rom_addr_offset + rom_addr_l2'length-1),
            scout   => sov(rom_addr_offset to rom_addr_offset + rom_addr_l2'length-1),
            din     => rom_addr_d,
            dout    => rom_addr_l2);
-----------------------------------------------------------------------
-- Scan
-----------------------------------------------------------------------
siv(0 TO scan_right) <=  sov(1 to scan_right) & scan_in;
scan_out  <=  sov(0);
END IUQ_UC_ROM;
