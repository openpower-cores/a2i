-- © IBM Corp. 2020
-- This softcore is licensed under and subject to the terms of the CC-BY 4.0
-- license (https://creativecommons.org/licenses/by/4.0/legalcode). 
-- Additional rights, including the right to physically implement a softcore 
-- that is compliant with the required sections of the Power ISA 
-- Specification, will be available at no cost via the OpenPOWER Foundation. 
-- This README will be updated with additional information when OpenPOWER's 
-- license is available.

			

library ieee,ibm,support,tri;
use ieee.std_logic_1164.all;
use ibm.std_ulogic_unsigned.all;
use ibm.std_ulogic_support.all;
use ibm.std_ulogic_function_support.all;
use support.power_logic_pkg.all;
use tri.tri_latches_pkg.all;

entity iuq_uc_rom is
  generic(ucode_width           : integer := 71;
          regmode               : integer := 6;
          expand_type           : integer := 2);
port(
     vdd                        : inout power_logic;
     gnd                        : inout power_logic;
     nclk                       : in clk_logic;
     pc_iu_func_sl_thold_0_b    : in std_ulogic;
     pc_iu_sg_0                 : in std_ulogic;
     forcee : in std_ulogic;
     d_mode                     : in std_ulogic;
     delay_lclkr                : in std_ulogic;
     mpw1_b                     : in std_ulogic;
     mpw2_b                     : in std_ulogic;
     scan_in                    : in std_ulogic;
     scan_out                   : out std_ulogic;

     rom_act                    : in std_ulogic;
     rom_addr                   : in std_ulogic_vector(0 to 9);
     rom_data                   : out std_ulogic_vector(0 to ucode_width-1)
);
-- synopsys translate_off
-- synopsys translate_on
end iuq_uc_rom;
ARCHITECTURE IUQ_UC_ROM
          OF IUQ_UC_ROM
          IS
SIGNAL ROM32_INSTR_PT                    : STD_ULOGIC_VECTOR(1 TO 893)  := 
(OTHERS=> 'U');
SIGNAL ROM64_INSTR_PT                    : STD_ULOGIC_VECTOR(1 TO 890)  := 
(OTHERS=> 'U');
SIGNAL count_src                         : STD_ULOGIC_VECTOR(0 TO 2)  := 
"UUU";
SIGNAL cr_bf2fxm                         : STD_ULOGIC  := 
'U';
SIGNAL ep                                : STD_ULOGIC  := 
'U';
SIGNAL extRT                             : STD_ULOGIC  := 
'U';
SIGNAL extS1                             : STD_ULOGIC  := 
'U';
SIGNAL extS2                             : STD_ULOGIC  := 
'U';
SIGNAL extS3                             : STD_ULOGIC  := 
'U';
SIGNAL loop_addr                         : STD_ULOGIC_VECTOR(0 TO 9)  := 
"UUUUUUUUUU";
SIGNAL loop_begin                        : STD_ULOGIC  := 
'U';
SIGNAL loop_end                          : STD_ULOGIC  := 
'U';
SIGNAL loop_init                         : STD_ULOGIC_VECTOR(0 TO 2)  := 
"UUU";
SIGNAL sel0_5                            : STD_ULOGIC  := 
'U';
SIGNAL sel11_15                          : STD_ULOGIC_VECTOR(0 TO 1)  := 
"UU";
SIGNAL sel16_20                          : STD_ULOGIC_VECTOR(0 TO 1)  := 
"UU";
SIGNAL sel21_25                          : STD_ULOGIC_VECTOR(0 TO 1)  := 
"UU";
SIGNAL sel26_30                          : STD_ULOGIC  := 
'U';
SIGNAL sel31                             : STD_ULOGIC  := 
'U';
SIGNAL sel6_10                           : STD_ULOGIC_VECTOR(0 TO 1)  := 
"UU";
SIGNAL skip_cond                         : STD_ULOGIC  := 
'U';
SIGNAL skip_zero                         : STD_ULOGIC  := 
'U';
SIGNAL template                          : STD_ULOGIC_VECTOR(0 TO 31)  := 
"UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU";
SIGNAL ucode_end                         : STD_ULOGIC  := 
'U';
SIGNAL ucode_end_early                   : STD_ULOGIC  := 
'U';
constant rom_addr_offset        : natural := 0;
constant scan_right             : natural := rom_addr_offset + 10 - 1;
signal rom_addr_d               : std_ulogic_vector(0 to 9);
signal rom_addr_l2              : std_ulogic_vector(0 to 9);
signal siv              : std_ulogic_vector(0 to scan_right);
signal sov              : std_ulogic_vector(0 to scan_right);
signal rom_unused       : std_ulogic;
-- synopsys translate_off
-- synopsys translate_on
  BEGIN 

c64: if (regmode = 6) generate
begin


ROM32_INSTR_PT  <=  (others => '0');
rom_unused  <=  or_reduce(ROM32_INSTR_PT);
MQQ1:ROM64_INSTR_PT(1) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100000000"));
MQQ2:ROM64_INSTR_PT(2) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000000"));
MQQ3:ROM64_INSTR_PT(3) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000000"));
MQQ4:ROM64_INSTR_PT(4) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000000"));
MQQ5:ROM64_INSTR_PT(5) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000000"));
MQQ6:ROM64_INSTR_PT(6) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110000000"));
MQQ7:ROM64_INSTR_PT(7) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000000"));
MQQ8:ROM64_INSTR_PT(8) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00100000"));
MQQ9:ROM64_INSTR_PT(9) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100000"));
MQQ10:ROM64_INSTR_PT(10) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100000"));
MQQ11:ROM64_INSTR_PT(11) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100000"));
MQQ12:ROM64_INSTR_PT(12) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000000"));
MQQ13:ROM64_INSTR_PT(13) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000000"));
MQQ14:ROM64_INSTR_PT(14) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010000"));
MQQ15:ROM64_INSTR_PT(15) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010000"));
MQQ16:ROM64_INSTR_PT(16) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101010000"));
MQQ17:ROM64_INSTR_PT(17) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000110000"));
MQQ18:ROM64_INSTR_PT(18) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010110000"));
MQQ19:ROM64_INSTR_PT(19) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0110000"));
MQQ20:ROM64_INSTR_PT(20) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110000"));
MQQ21:ROM64_INSTR_PT(21) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110000"));
MQQ22:ROM64_INSTR_PT(22) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110000"));
MQQ23:ROM64_INSTR_PT(23) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010000"));
MQQ24:ROM64_INSTR_PT(24) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110000"));
MQQ25:ROM64_INSTR_PT(25) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ26:ROM64_INSTR_PT(26) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000000"));
MQQ27:ROM64_INSTR_PT(27) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100000"));
MQQ28:ROM64_INSTR_PT(28) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010000"));
MQQ29:ROM64_INSTR_PT(29) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110000"));
MQQ30:ROM64_INSTR_PT(30) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ31:ROM64_INSTR_PT(31) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110000"));
MQQ32:ROM64_INSTR_PT(32) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0010000"));
MQQ33:ROM64_INSTR_PT(33) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010000"));
MQQ34:ROM64_INSTR_PT(34) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010000"));
MQQ35:ROM64_INSTR_PT(35) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110000"));
MQQ36:ROM64_INSTR_PT(36) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001000"));
MQQ37:ROM64_INSTR_PT(37) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101001000"));
MQQ38:ROM64_INSTR_PT(38) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110001000"));
MQQ39:ROM64_INSTR_PT(39) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001000"));
MQQ40:ROM64_INSTR_PT(40) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101000"));
MQQ41:ROM64_INSTR_PT(41) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001101000"));
MQQ42:ROM64_INSTR_PT(42) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101000"));
MQQ43:ROM64_INSTR_PT(43) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101000"));
MQQ44:ROM64_INSTR_PT(44) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101000"));
MQQ45:ROM64_INSTR_PT(45) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111101000"));
MQQ46:ROM64_INSTR_PT(46) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001000"));
MQQ47:ROM64_INSTR_PT(47) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101000"));
MQQ48:ROM64_INSTR_PT(48) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001011000"));
MQQ49:ROM64_INSTR_PT(49) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011011000"));
MQQ50:ROM64_INSTR_PT(50) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011000"));
MQQ51:ROM64_INSTR_PT(51) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111000"));
MQQ52:ROM64_INSTR_PT(52) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111000"));
MQQ53:ROM64_INSTR_PT(53) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111000"));
MQQ54:ROM64_INSTR_PT(54) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011000"));
MQQ55:ROM64_INSTR_PT(55) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111000"));
MQQ56:ROM64_INSTR_PT(56) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111000"));
MQQ57:ROM64_INSTR_PT(57) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111000"));
MQQ58:ROM64_INSTR_PT(58) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001000"));
MQQ59:ROM64_INSTR_PT(59) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011000"));
MQQ60:ROM64_INSTR_PT(60) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011000"));
MQQ61:ROM64_INSTR_PT(61) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100111000"));
MQQ62:ROM64_INSTR_PT(62) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111000"));
MQQ63:ROM64_INSTR_PT(63) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000000"));
MQQ64:ROM64_INSTR_PT(64) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000000"));
MQQ65:ROM64_INSTR_PT(65) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000000"));
MQQ66:ROM64_INSTR_PT(66) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010000"));
MQQ67:ROM64_INSTR_PT(67) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ68:ROM64_INSTR_PT(68) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100000"));
MQQ69:ROM64_INSTR_PT(69) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010000"));
MQQ70:ROM64_INSTR_PT(70) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001000"));
MQQ71:ROM64_INSTR_PT(71) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011000"));
MQQ72:ROM64_INSTR_PT(72) <=
    Eq(( ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000"));
MQQ73:ROM64_INSTR_PT(73) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100000100"));
MQQ74:ROM64_INSTR_PT(74) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000100"));
MQQ75:ROM64_INSTR_PT(75) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000100"));
MQQ76:ROM64_INSTR_PT(76) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000100"));
MQQ77:ROM64_INSTR_PT(77) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000100"));
MQQ78:ROM64_INSTR_PT(78) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000100"));
MQQ79:ROM64_INSTR_PT(79) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000100"));
MQQ80:ROM64_INSTR_PT(80) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100100100"));
MQQ81:ROM64_INSTR_PT(81) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100100"));
MQQ82:ROM64_INSTR_PT(82) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100100"));
MQQ83:ROM64_INSTR_PT(83) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100100"));
MQQ84:ROM64_INSTR_PT(84) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11100100"));
MQQ85:ROM64_INSTR_PT(85) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100100"));
MQQ86:ROM64_INSTR_PT(86) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000100"));
MQQ87:ROM64_INSTR_PT(87) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000100"));
MQQ88:ROM64_INSTR_PT(88) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100100"));
MQQ89:ROM64_INSTR_PT(89) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100010100"));
MQQ90:ROM64_INSTR_PT(90) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110010100"));
MQQ91:ROM64_INSTR_PT(91) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010100"));
MQQ92:ROM64_INSTR_PT(92) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010100"));
MQQ93:ROM64_INSTR_PT(93) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010100"));
MQQ94:ROM64_INSTR_PT(94) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010100"));
MQQ95:ROM64_INSTR_PT(95) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000110100"));
MQQ96:ROM64_INSTR_PT(96) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010110100"));
MQQ97:ROM64_INSTR_PT(97) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110100"));
MQQ98:ROM64_INSTR_PT(98) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110100"));
MQQ99:ROM64_INSTR_PT(99) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110100"));
MQQ100:ROM64_INSTR_PT(100) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110100"));
MQQ101:ROM64_INSTR_PT(101) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110100"));
MQQ102:ROM64_INSTR_PT(102) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000100"));
MQQ103:ROM64_INSTR_PT(103) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010100"));
MQQ104:ROM64_INSTR_PT(104) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110100"));
MQQ105:ROM64_INSTR_PT(105) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010100"));
MQQ106:ROM64_INSTR_PT(106) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100001100"));
MQQ107:ROM64_INSTR_PT(107) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001001100"));
MQQ108:ROM64_INSTR_PT(108) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001001100"));
MQQ109:ROM64_INSTR_PT(109) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001100"));
MQQ110:ROM64_INSTR_PT(110) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001100"));
MQQ111:ROM64_INSTR_PT(111) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001100"));
MQQ112:ROM64_INSTR_PT(112) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101100"));
MQQ113:ROM64_INSTR_PT(113) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100101100"));
MQQ114:ROM64_INSTR_PT(114) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010101100"));
MQQ115:ROM64_INSTR_PT(115) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101100"));
MQQ116:ROM64_INSTR_PT(116) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101100"));
MQQ117:ROM64_INSTR_PT(117) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ118:ROM64_INSTR_PT(118) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ119:ROM64_INSTR_PT(119) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011100"));
MQQ120:ROM64_INSTR_PT(120) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011100"));
MQQ121:ROM64_INSTR_PT(121) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011011100"));
MQQ122:ROM64_INSTR_PT(122) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ123:ROM64_INSTR_PT(123) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100111100"));
MQQ124:ROM64_INSTR_PT(124) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111100"));
MQQ125:ROM64_INSTR_PT(125) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ126:ROM64_INSTR_PT(126) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ127:ROM64_INSTR_PT(127) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011100"));
MQQ128:ROM64_INSTR_PT(128) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011100"));
MQQ129:ROM64_INSTR_PT(129) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111100"));
MQQ130:ROM64_INSTR_PT(130) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ131:ROM64_INSTR_PT(131) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011100"));
MQQ132:ROM64_INSTR_PT(132) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ133:ROM64_INSTR_PT(133) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001100"));
MQQ134:ROM64_INSTR_PT(134) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101100"));
MQQ135:ROM64_INSTR_PT(135) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ136:ROM64_INSTR_PT(136) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111100"));
MQQ137:ROM64_INSTR_PT(137) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111100"));
MQQ138:ROM64_INSTR_PT(138) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0100100"));
MQQ139:ROM64_INSTR_PT(139) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010100"));
MQQ140:ROM64_INSTR_PT(140) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010100"));
MQQ141:ROM64_INSTR_PT(141) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001100"));
MQQ142:ROM64_INSTR_PT(142) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001100"));
MQQ143:ROM64_INSTR_PT(143) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ144:ROM64_INSTR_PT(144) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111100"));
MQQ145:ROM64_INSTR_PT(145) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ146:ROM64_INSTR_PT(146) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001100"));
MQQ147:ROM64_INSTR_PT(147) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000000"));
MQQ148:ROM64_INSTR_PT(148) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010000"));
MQQ149:ROM64_INSTR_PT(149) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010000"));
MQQ150:ROM64_INSTR_PT(150) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001000"));
MQQ151:ROM64_INSTR_PT(151) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001000"));
MQQ152:ROM64_INSTR_PT(152) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1000"));
MQQ153:ROM64_INSTR_PT(153) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000100"));
MQQ154:ROM64_INSTR_PT(154) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000100"));
MQQ155:ROM64_INSTR_PT(155) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100100"));
MQQ156:ROM64_INSTR_PT(156) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("00100"));
MQQ157:ROM64_INSTR_PT(157) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ158:ROM64_INSTR_PT(158) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ159:ROM64_INSTR_PT(159) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111100"));
MQQ160:ROM64_INSTR_PT(160) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011100"));
MQQ161:ROM64_INSTR_PT(161) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011100"));
MQQ162:ROM64_INSTR_PT(162) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111100"));
MQQ163:ROM64_INSTR_PT(163) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("01000"));
MQQ164:ROM64_INSTR_PT(164) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000100"));
MQQ165:ROM64_INSTR_PT(165) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("10100"));
MQQ166:ROM64_INSTR_PT(166) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ167:ROM64_INSTR_PT(167) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("01100"));
MQQ168:ROM64_INSTR_PT(168) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100000010"));
MQQ169:ROM64_INSTR_PT(169) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000010"));
MQQ170:ROM64_INSTR_PT(170) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000010"));
MQQ171:ROM64_INSTR_PT(171) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000010"));
MQQ172:ROM64_INSTR_PT(172) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000010"));
MQQ173:ROM64_INSTR_PT(173) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100010"));
MQQ174:ROM64_INSTR_PT(174) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100010"));
MQQ175:ROM64_INSTR_PT(175) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100010"));
MQQ176:ROM64_INSTR_PT(176) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000010"));
MQQ177:ROM64_INSTR_PT(177) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ178:ROM64_INSTR_PT(178) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("000010"));
MQQ179:ROM64_INSTR_PT(179) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010010"));
MQQ180:ROM64_INSTR_PT(180) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001110010"));
MQQ181:ROM64_INSTR_PT(181) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110010"));
MQQ182:ROM64_INSTR_PT(182) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110010"));
MQQ183:ROM64_INSTR_PT(183) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110010"));
MQQ184:ROM64_INSTR_PT(184) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010010"));
MQQ185:ROM64_INSTR_PT(185) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010010"));
MQQ186:ROM64_INSTR_PT(186) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110010"));
MQQ187:ROM64_INSTR_PT(187) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110010"));
MQQ188:ROM64_INSTR_PT(188) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ189:ROM64_INSTR_PT(189) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000010"));
MQQ190:ROM64_INSTR_PT(190) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000010"));
MQQ191:ROM64_INSTR_PT(191) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100010"));
MQQ192:ROM64_INSTR_PT(192) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ193:ROM64_INSTR_PT(193) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110010"));
MQQ194:ROM64_INSTR_PT(194) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110010"));
MQQ195:ROM64_INSTR_PT(195) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110010"));
MQQ196:ROM64_INSTR_PT(196) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ197:ROM64_INSTR_PT(197) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110010"));
MQQ198:ROM64_INSTR_PT(198) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ199:ROM64_INSTR_PT(199) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001010"));
MQQ200:ROM64_INSTR_PT(200) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101001010"));
MQQ201:ROM64_INSTR_PT(201) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001001010"));
MQQ202:ROM64_INSTR_PT(202) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001010"));
MQQ203:ROM64_INSTR_PT(203) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001010"));
MQQ204:ROM64_INSTR_PT(204) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001010"));
MQQ205:ROM64_INSTR_PT(205) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101010"));
MQQ206:ROM64_INSTR_PT(206) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101010"));
MQQ207:ROM64_INSTR_PT(207) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101010"));
MQQ208:ROM64_INSTR_PT(208) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101010"));
MQQ209:ROM64_INSTR_PT(209) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101010"));
MQQ210:ROM64_INSTR_PT(210) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001010"));
MQQ211:ROM64_INSTR_PT(211) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011010"));
MQQ212:ROM64_INSTR_PT(212) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ213:ROM64_INSTR_PT(213) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011010"));
MQQ214:ROM64_INSTR_PT(214) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011011010"));
MQQ215:ROM64_INSTR_PT(215) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111010"));
MQQ216:ROM64_INSTR_PT(216) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011111010"));
MQQ217:ROM64_INSTR_PT(217) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111010"));
MQQ218:ROM64_INSTR_PT(218) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111010"));
MQQ219:ROM64_INSTR_PT(219) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011010"));
MQQ220:ROM64_INSTR_PT(220) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011010"));
MQQ221:ROM64_INSTR_PT(221) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100111010"));
MQQ222:ROM64_INSTR_PT(222) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111010"));
MQQ223:ROM64_INSTR_PT(223) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111010"));
MQQ224:ROM64_INSTR_PT(224) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101010"));
MQQ225:ROM64_INSTR_PT(225) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011010"));
MQQ226:ROM64_INSTR_PT(226) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ227:ROM64_INSTR_PT(227) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011010"));
MQQ228:ROM64_INSTR_PT(228) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100010"));
MQQ229:ROM64_INSTR_PT(229) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100010"));
MQQ230:ROM64_INSTR_PT(230) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010010"));
MQQ231:ROM64_INSTR_PT(231) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ232:ROM64_INSTR_PT(232) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001010"));
MQQ233:ROM64_INSTR_PT(233) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101010"));
MQQ234:ROM64_INSTR_PT(234) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011010"));
MQQ235:ROM64_INSTR_PT(235) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011010"));
MQQ236:ROM64_INSTR_PT(236) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100000110"));
MQQ237:ROM64_INSTR_PT(237) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110000110"));
MQQ238:ROM64_INSTR_PT(238) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000110"));
MQQ239:ROM64_INSTR_PT(239) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000110"));
MQQ240:ROM64_INSTR_PT(240) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000110"));
MQQ241:ROM64_INSTR_PT(241) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000110"));
MQQ242:ROM64_INSTR_PT(242) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111000110"));
MQQ243:ROM64_INSTR_PT(243) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000110"));
MQQ244:ROM64_INSTR_PT(244) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000110"));
MQQ245:ROM64_INSTR_PT(245) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000100110"));
MQQ246:ROM64_INSTR_PT(246) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100110"));
MQQ247:ROM64_INSTR_PT(247) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001100110"));
MQQ248:ROM64_INSTR_PT(248) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000110"));
MQQ249:ROM64_INSTR_PT(249) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000110"));
MQQ250:ROM64_INSTR_PT(250) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000110"));
MQQ251:ROM64_INSTR_PT(251) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100110"));
MQQ252:ROM64_INSTR_PT(252) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110010110"));
MQQ253:ROM64_INSTR_PT(253) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010110"));
MQQ254:ROM64_INSTR_PT(254) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010110"));
MQQ255:ROM64_INSTR_PT(255) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110110"));
MQQ256:ROM64_INSTR_PT(256) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110110"));
MQQ257:ROM64_INSTR_PT(257) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110110"));
MQQ258:ROM64_INSTR_PT(258) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110110"));
MQQ259:ROM64_INSTR_PT(259) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100110110"));
MQQ260:ROM64_INSTR_PT(260) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110110"));
MQQ261:ROM64_INSTR_PT(261) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110110"));
MQQ262:ROM64_INSTR_PT(262) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100110"));
MQQ263:ROM64_INSTR_PT(263) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100110110"));
MQQ264:ROM64_INSTR_PT(264) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110110"));
MQQ265:ROM64_INSTR_PT(265) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100001110"));
MQQ266:ROM64_INSTR_PT(266) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001110"));
MQQ267:ROM64_INSTR_PT(267) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110001110"));
MQQ268:ROM64_INSTR_PT(268) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001110"));
MQQ269:ROM64_INSTR_PT(269) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001110"));
MQQ270:ROM64_INSTR_PT(270) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000101110"));
MQQ271:ROM64_INSTR_PT(271) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100101110"));
MQQ272:ROM64_INSTR_PT(272) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101110"));
MQQ273:ROM64_INSTR_PT(273) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101110"));
MQQ274:ROM64_INSTR_PT(274) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101110"));
MQQ275:ROM64_INSTR_PT(275) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101110"));
MQQ276:ROM64_INSTR_PT(276) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101110"));
MQQ277:ROM64_INSTR_PT(277) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011110"));
MQQ278:ROM64_INSTR_PT(278) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011110"));
MQQ279:ROM64_INSTR_PT(279) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ280:ROM64_INSTR_PT(280) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111110"));
MQQ281:ROM64_INSTR_PT(281) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111110"));
MQQ282:ROM64_INSTR_PT(282) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111110"));
MQQ283:ROM64_INSTR_PT(283) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011110"));
MQQ284:ROM64_INSTR_PT(284) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011110"));
MQQ285:ROM64_INSTR_PT(285) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ286:ROM64_INSTR_PT(286) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111110"));
MQQ287:ROM64_INSTR_PT(287) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111110"));
MQQ288:ROM64_INSTR_PT(288) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111110"));
MQQ289:ROM64_INSTR_PT(289) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111110"));
MQQ290:ROM64_INSTR_PT(290) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ291:ROM64_INSTR_PT(291) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111110"));
MQQ292:ROM64_INSTR_PT(292) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111110"));
MQQ293:ROM64_INSTR_PT(293) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ294:ROM64_INSTR_PT(294) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110110"));
MQQ295:ROM64_INSTR_PT(295) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100110"));
MQQ296:ROM64_INSTR_PT(296) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001110"));
MQQ297:ROM64_INSTR_PT(297) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ298:ROM64_INSTR_PT(298) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111110"));
MQQ299:ROM64_INSTR_PT(299) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011110"));
MQQ300:ROM64_INSTR_PT(300) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ301:ROM64_INSTR_PT(301) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101110"));
MQQ302:ROM64_INSTR_PT(302) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101110"));
MQQ303:ROM64_INSTR_PT(303) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000010"));
MQQ304:ROM64_INSTR_PT(304) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011010"));
MQQ305:ROM64_INSTR_PT(305) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ306:ROM64_INSTR_PT(306) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ307:ROM64_INSTR_PT(307) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101010"));
MQQ308:ROM64_INSTR_PT(308) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000110"));
MQQ309:ROM64_INSTR_PT(309) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000110"));
MQQ310:ROM64_INSTR_PT(310) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010110"));
MQQ311:ROM64_INSTR_PT(311) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110110"));
MQQ312:ROM64_INSTR_PT(312) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001110"));
MQQ313:ROM64_INSTR_PT(313) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001110"));
MQQ314:ROM64_INSTR_PT(314) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111110"));
MQQ315:ROM64_INSTR_PT(315) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ316:ROM64_INSTR_PT(316) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010110"));
MQQ317:ROM64_INSTR_PT(317) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010010"));
MQQ318:ROM64_INSTR_PT(318) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("01010"));
MQQ319:ROM64_INSTR_PT(319) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ320:ROM64_INSTR_PT(320) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0000010"));
MQQ321:ROM64_INSTR_PT(321) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000000"));
MQQ322:ROM64_INSTR_PT(322) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010000"));
MQQ323:ROM64_INSTR_PT(323) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000000"));
MQQ324:ROM64_INSTR_PT(324) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101000"));
MQQ325:ROM64_INSTR_PT(325) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101000"));
MQQ326:ROM64_INSTR_PT(326) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101000"));
MQQ327:ROM64_INSTR_PT(327) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100000"));
MQQ328:ROM64_INSTR_PT(328) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011000"));
MQQ329:ROM64_INSTR_PT(329) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0000100"));
MQQ330:ROM64_INSTR_PT(330) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000100"));
MQQ331:ROM64_INSTR_PT(331) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000100"));
MQQ332:ROM64_INSTR_PT(332) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000100"));
MQQ333:ROM64_INSTR_PT(333) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001100"));
MQQ334:ROM64_INSTR_PT(334) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00101100"));
MQQ335:ROM64_INSTR_PT(335) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011100"));
MQQ336:ROM64_INSTR_PT(336) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000000"));
MQQ337:ROM64_INSTR_PT(337) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ338:ROM64_INSTR_PT(338) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000010"));
MQQ339:ROM64_INSTR_PT(339) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ340:ROM64_INSTR_PT(340) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010010"));
MQQ341:ROM64_INSTR_PT(341) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ342:ROM64_INSTR_PT(342) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ343:ROM64_INSTR_PT(343) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001010"));
MQQ344:ROM64_INSTR_PT(344) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001010"));
MQQ345:ROM64_INSTR_PT(345) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100110"));
MQQ346:ROM64_INSTR_PT(346) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ347:ROM64_INSTR_PT(347) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ348:ROM64_INSTR_PT(348) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ349:ROM64_INSTR_PT(349) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101110"));
MQQ350:ROM64_INSTR_PT(350) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ351:ROM64_INSTR_PT(351) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101010"));
MQQ352:ROM64_INSTR_PT(352) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101110"));
MQQ353:ROM64_INSTR_PT(353) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011110"));
MQQ354:ROM64_INSTR_PT(354) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000000"));
MQQ355:ROM64_INSTR_PT(355) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ356:ROM64_INSTR_PT(356) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000010"));
MQQ357:ROM64_INSTR_PT(357) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100010"));
MQQ358:ROM64_INSTR_PT(358) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110110"));
MQQ359:ROM64_INSTR_PT(359) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011110"));
MQQ360:ROM64_INSTR_PT(360) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100010"));
MQQ361:ROM64_INSTR_PT(361) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100000001"));
MQQ362:ROM64_INSTR_PT(362) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000001"));
MQQ363:ROM64_INSTR_PT(363) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000001"));
MQQ364:ROM64_INSTR_PT(364) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110000001"));
MQQ365:ROM64_INSTR_PT(365) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000001"));
MQQ366:ROM64_INSTR_PT(366) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100001"));
MQQ367:ROM64_INSTR_PT(367) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11100001"));
MQQ368:ROM64_INSTR_PT(368) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000001"));
MQQ369:ROM64_INSTR_PT(369) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ370:ROM64_INSTR_PT(370) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010001"));
MQQ371:ROM64_INSTR_PT(371) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010001"));
MQQ372:ROM64_INSTR_PT(372) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010001"));
MQQ373:ROM64_INSTR_PT(373) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110001"));
MQQ374:ROM64_INSTR_PT(374) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010110001"));
MQQ375:ROM64_INSTR_PT(375) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001110001"));
MQQ376:ROM64_INSTR_PT(376) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00110001"));
MQQ377:ROM64_INSTR_PT(377) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110001"));
MQQ378:ROM64_INSTR_PT(378) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110001"));
MQQ379:ROM64_INSTR_PT(379) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110001"));
MQQ380:ROM64_INSTR_PT(380) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110001"));
MQQ381:ROM64_INSTR_PT(381) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110001"));
MQQ382:ROM64_INSTR_PT(382) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110001"));
MQQ383:ROM64_INSTR_PT(383) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ384:ROM64_INSTR_PT(384) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100001"));
MQQ385:ROM64_INSTR_PT(385) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100110001"));
MQQ386:ROM64_INSTR_PT(386) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110001"));
MQQ387:ROM64_INSTR_PT(387) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010001"));
MQQ388:ROM64_INSTR_PT(388) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001001"));
MQQ389:ROM64_INSTR_PT(389) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111001001"));
MQQ390:ROM64_INSTR_PT(390) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001001"));
MQQ391:ROM64_INSTR_PT(391) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001001"));
MQQ392:ROM64_INSTR_PT(392) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101001"));
MQQ393:ROM64_INSTR_PT(393) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00101001"));
MQQ394:ROM64_INSTR_PT(394) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101001"));
MQQ395:ROM64_INSTR_PT(395) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001101001"));
MQQ396:ROM64_INSTR_PT(396) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101001"));
MQQ397:ROM64_INSTR_PT(397) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101001"));
MQQ398:ROM64_INSTR_PT(398) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111101001"));
MQQ399:ROM64_INSTR_PT(399) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001001"));
MQQ400:ROM64_INSTR_PT(400) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("001001"));
MQQ401:ROM64_INSTR_PT(401) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011001"));
MQQ402:ROM64_INSTR_PT(402) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001011001"));
MQQ403:ROM64_INSTR_PT(403) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011111001"));
MQQ404:ROM64_INSTR_PT(404) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111001"));
MQQ405:ROM64_INSTR_PT(405) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011001"));
MQQ406:ROM64_INSTR_PT(406) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011001"));
MQQ407:ROM64_INSTR_PT(407) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011001"));
MQQ408:ROM64_INSTR_PT(408) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111001"));
MQQ409:ROM64_INSTR_PT(409) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111001"));
MQQ410:ROM64_INSTR_PT(410) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111001"));
MQQ411:ROM64_INSTR_PT(411) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011001"));
MQQ412:ROM64_INSTR_PT(412) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111001"));
MQQ413:ROM64_INSTR_PT(413) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111001"));
MQQ414:ROM64_INSTR_PT(414) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000001"));
MQQ415:ROM64_INSTR_PT(415) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ416:ROM64_INSTR_PT(416) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100001"));
MQQ417:ROM64_INSTR_PT(417) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010001"));
MQQ418:ROM64_INSTR_PT(418) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010001"));
MQQ419:ROM64_INSTR_PT(419) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101001"));
MQQ420:ROM64_INSTR_PT(420) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011001"));
MQQ421:ROM64_INSTR_PT(421) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011001"));
MQQ422:ROM64_INSTR_PT(422) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100000101"));
MQQ423:ROM64_INSTR_PT(423) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000101"));
MQQ424:ROM64_INSTR_PT(424) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000101"));
MQQ425:ROM64_INSTR_PT(425) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000101"));
MQQ426:ROM64_INSTR_PT(426) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000101"));
MQQ427:ROM64_INSTR_PT(427) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000101"));
MQQ428:ROM64_INSTR_PT(428) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000101"));
MQQ429:ROM64_INSTR_PT(429) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100100101"));
MQQ430:ROM64_INSTR_PT(430) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100101"));
MQQ431:ROM64_INSTR_PT(431) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100101"));
MQQ432:ROM64_INSTR_PT(432) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100101"));
MQQ433:ROM64_INSTR_PT(433) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100101"));
MQQ434:ROM64_INSTR_PT(434) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100101"));
MQQ435:ROM64_INSTR_PT(435) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11100101"));
MQQ436:ROM64_INSTR_PT(436) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100101"));
MQQ437:ROM64_INSTR_PT(437) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110010101"));
MQQ438:ROM64_INSTR_PT(438) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010101"));
MQQ439:ROM64_INSTR_PT(439) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101010101"));
MQQ440:ROM64_INSTR_PT(440) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010101"));
MQQ441:ROM64_INSTR_PT(441) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000110101"));
MQQ442:ROM64_INSTR_PT(442) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110101"));
MQQ443:ROM64_INSTR_PT(443) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110101"));
MQQ444:ROM64_INSTR_PT(444) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110101"));
MQQ445:ROM64_INSTR_PT(445) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110101"));
MQQ446:ROM64_INSTR_PT(446) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000101"));
MQQ447:ROM64_INSTR_PT(447) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100101"));
MQQ448:ROM64_INSTR_PT(448) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110101"));
MQQ449:ROM64_INSTR_PT(449) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110101"));
MQQ450:ROM64_INSTR_PT(450) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010101"));
MQQ451:ROM64_INSTR_PT(451) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100001101"));
MQQ452:ROM64_INSTR_PT(452) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110001101"));
MQQ453:ROM64_INSTR_PT(453) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001001101"));
MQQ454:ROM64_INSTR_PT(454) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001101"));
MQQ455:ROM64_INSTR_PT(455) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010101101"));
MQQ456:ROM64_INSTR_PT(456) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101101"));
MQQ457:ROM64_INSTR_PT(457) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101101"));
MQQ458:ROM64_INSTR_PT(458) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101101"));
MQQ459:ROM64_INSTR_PT(459) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001101"));
MQQ460:ROM64_INSTR_PT(460) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101101"));
MQQ461:ROM64_INSTR_PT(461) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011101"));
MQQ462:ROM64_INSTR_PT(462) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011101"));
MQQ463:ROM64_INSTR_PT(463) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111101"));
MQQ464:ROM64_INSTR_PT(464) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111101"));
MQQ465:ROM64_INSTR_PT(465) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011101"));
MQQ466:ROM64_INSTR_PT(466) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011101"));
MQQ467:ROM64_INSTR_PT(467) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111101"));
MQQ468:ROM64_INSTR_PT(468) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100111101"));
MQQ469:ROM64_INSTR_PT(469) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111101"));
MQQ470:ROM64_INSTR_PT(470) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111101"));
MQQ471:ROM64_INSTR_PT(471) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001101"));
MQQ472:ROM64_INSTR_PT(472) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100101"));
MQQ473:ROM64_INSTR_PT(473) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010101"));
MQQ474:ROM64_INSTR_PT(474) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110101"));
MQQ475:ROM64_INSTR_PT(475) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010101"));
MQQ476:ROM64_INSTR_PT(476) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010101"));
MQQ477:ROM64_INSTR_PT(477) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001101"));
MQQ478:ROM64_INSTR_PT(478) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001101"));
MQQ479:ROM64_INSTR_PT(479) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001101"));
MQQ480:ROM64_INSTR_PT(480) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011101"));
MQQ481:ROM64_INSTR_PT(481) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111101"));
MQQ482:ROM64_INSTR_PT(482) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ483:ROM64_INSTR_PT(483) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010001"));
MQQ484:ROM64_INSTR_PT(484) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110001"));
MQQ485:ROM64_INSTR_PT(485) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001001"));
MQQ486:ROM64_INSTR_PT(486) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001001"));
MQQ487:ROM64_INSTR_PT(487) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101001"));
MQQ488:ROM64_INSTR_PT(488) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011001"));
MQQ489:ROM64_INSTR_PT(489) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111001"));
MQQ490:ROM64_INSTR_PT(490) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111001"));
MQQ491:ROM64_INSTR_PT(491) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000101"));
MQQ492:ROM64_INSTR_PT(492) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100101"));
MQQ493:ROM64_INSTR_PT(493) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100101"));
MQQ494:ROM64_INSTR_PT(494) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100101"));
MQQ495:ROM64_INSTR_PT(495) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111101"));
MQQ496:ROM64_INSTR_PT(496) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011101"));
MQQ497:ROM64_INSTR_PT(497) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111101"));
MQQ498:ROM64_INSTR_PT(498) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101101"));
MQQ499:ROM64_INSTR_PT(499) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001101"));
MQQ500:ROM64_INSTR_PT(500) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0000001"));
MQQ501:ROM64_INSTR_PT(501) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("001101"));
MQQ502:ROM64_INSTR_PT(502) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001"));
MQQ503:ROM64_INSTR_PT(503) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100000011"));
MQQ504:ROM64_INSTR_PT(504) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000011"));
MQQ505:ROM64_INSTR_PT(505) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000011"));
MQQ506:ROM64_INSTR_PT(506) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000011"));
MQQ507:ROM64_INSTR_PT(507) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000011"));
MQQ508:ROM64_INSTR_PT(508) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010100011"));
MQQ509:ROM64_INSTR_PT(509) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100011"));
MQQ510:ROM64_INSTR_PT(510) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100011"));
MQQ511:ROM64_INSTR_PT(511) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000011"));
MQQ512:ROM64_INSTR_PT(512) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100011"));
MQQ513:ROM64_INSTR_PT(513) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000011"));
MQQ514:ROM64_INSTR_PT(514) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010011"));
MQQ515:ROM64_INSTR_PT(515) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010011"));
MQQ516:ROM64_INSTR_PT(516) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010011"));
MQQ517:ROM64_INSTR_PT(517) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010011"));
MQQ518:ROM64_INSTR_PT(518) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010011"));
MQQ519:ROM64_INSTR_PT(519) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001110011"));
MQQ520:ROM64_INSTR_PT(520) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110011"));
MQQ521:ROM64_INSTR_PT(521) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110011"));
MQQ522:ROM64_INSTR_PT(522) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110011"));
MQQ523:ROM64_INSTR_PT(523) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110011"));
MQQ524:ROM64_INSTR_PT(524) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000011"));
MQQ525:ROM64_INSTR_PT(525) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100011"));
MQQ526:ROM64_INSTR_PT(526) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100011"));
MQQ527:ROM64_INSTR_PT(527) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010011"));
MQQ528:ROM64_INSTR_PT(528) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110011"));
MQQ529:ROM64_INSTR_PT(529) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010011"));
MQQ530:ROM64_INSTR_PT(530) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001011"));
MQQ531:ROM64_INSTR_PT(531) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101001011"));
MQQ532:ROM64_INSTR_PT(532) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001001011"));
MQQ533:ROM64_INSTR_PT(533) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111001011"));
MQQ534:ROM64_INSTR_PT(534) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000101011"));
MQQ535:ROM64_INSTR_PT(535) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101011"));
MQQ536:ROM64_INSTR_PT(536) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001101011"));
MQQ537:ROM64_INSTR_PT(537) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101011"));
MQQ538:ROM64_INSTR_PT(538) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101011"));
MQQ539:ROM64_INSTR_PT(539) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001011"));
MQQ540:ROM64_INSTR_PT(540) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101011"));
MQQ541:ROM64_INSTR_PT(541) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011011"));
MQQ542:ROM64_INSTR_PT(542) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ543:ROM64_INSTR_PT(543) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011011"));
MQQ544:ROM64_INSTR_PT(544) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111011"));
MQQ545:ROM64_INSTR_PT(545) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011011"));
MQQ546:ROM64_INSTR_PT(546) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011011"));
MQQ547:ROM64_INSTR_PT(547) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ548:ROM64_INSTR_PT(548) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111011"));
MQQ549:ROM64_INSTR_PT(549) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101011"));
MQQ550:ROM64_INSTR_PT(550) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011011"));
MQQ551:ROM64_INSTR_PT(551) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ552:ROM64_INSTR_PT(552) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100011"));
MQQ553:ROM64_INSTR_PT(553) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100011"));
MQQ554:ROM64_INSTR_PT(554) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010011"));
MQQ555:ROM64_INSTR_PT(555) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110011"));
MQQ556:ROM64_INSTR_PT(556) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001011"));
MQQ557:ROM64_INSTR_PT(557) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101011"));
MQQ558:ROM64_INSTR_PT(558) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011011"));
MQQ559:ROM64_INSTR_PT(559) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011011"));
MQQ560:ROM64_INSTR_PT(560) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111011"));
MQQ561:ROM64_INSTR_PT(561) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101011"));
MQQ562:ROM64_INSTR_PT(562) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011011"));
MQQ563:ROM64_INSTR_PT(563) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111011"));
MQQ564:ROM64_INSTR_PT(564) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111011"));
MQQ565:ROM64_INSTR_PT(565) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ566:ROM64_INSTR_PT(566) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000111"));
MQQ567:ROM64_INSTR_PT(567) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000111"));
MQQ568:ROM64_INSTR_PT(568) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110000111"));
MQQ569:ROM64_INSTR_PT(569) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000111"));
MQQ570:ROM64_INSTR_PT(570) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000111"));
MQQ571:ROM64_INSTR_PT(571) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000111"));
MQQ572:ROM64_INSTR_PT(572) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010100111"));
MQQ573:ROM64_INSTR_PT(573) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100111"));
MQQ574:ROM64_INSTR_PT(574) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100111"));
MQQ575:ROM64_INSTR_PT(575) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100111"));
MQQ576:ROM64_INSTR_PT(576) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100111"));
MQQ577:ROM64_INSTR_PT(577) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100111"));
MQQ578:ROM64_INSTR_PT(578) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000111"));
MQQ579:ROM64_INSTR_PT(579) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010111"));
MQQ580:ROM64_INSTR_PT(580) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010111"));
MQQ581:ROM64_INSTR_PT(581) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001010111"));
MQQ582:ROM64_INSTR_PT(582) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010111"));
MQQ583:ROM64_INSTR_PT(583) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110111"));
MQQ584:ROM64_INSTR_PT(584) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010111"));
MQQ585:ROM64_INSTR_PT(585) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000111"));
MQQ586:ROM64_INSTR_PT(586) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100111"));
MQQ587:ROM64_INSTR_PT(587) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010111"));
MQQ588:ROM64_INSTR_PT(588) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001111"));
MQQ589:ROM64_INSTR_PT(589) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100001111"));
MQQ590:ROM64_INSTR_PT(590) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001111"));
MQQ591:ROM64_INSTR_PT(591) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001111"));
MQQ592:ROM64_INSTR_PT(592) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001111"));
MQQ593:ROM64_INSTR_PT(593) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001111"));
MQQ594:ROM64_INSTR_PT(594) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001111"));
MQQ595:ROM64_INSTR_PT(595) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000101111"));
MQQ596:ROM64_INSTR_PT(596) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010101111"));
MQQ597:ROM64_INSTR_PT(597) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001101111"));
MQQ598:ROM64_INSTR_PT(598) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101111"));
MQQ599:ROM64_INSTR_PT(599) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101111"));
MQQ600:ROM64_INSTR_PT(600) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101111"));
MQQ601:ROM64_INSTR_PT(601) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011111"));
MQQ602:ROM64_INSTR_PT(602) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011111"));
MQQ603:ROM64_INSTR_PT(603) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001011111"));
MQQ604:ROM64_INSTR_PT(604) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111111"));
MQQ605:ROM64_INSTR_PT(605) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111111"));
MQQ606:ROM64_INSTR_PT(606) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111111"));
MQQ607:ROM64_INSTR_PT(607) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ608:ROM64_INSTR_PT(608) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011111"));
MQQ609:ROM64_INSTR_PT(609) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ610:ROM64_INSTR_PT(610) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111111"));
MQQ611:ROM64_INSTR_PT(611) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111111"));
MQQ612:ROM64_INSTR_PT(612) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111111"));
MQQ613:ROM64_INSTR_PT(613) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101111"));
MQQ614:ROM64_INSTR_PT(614) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ615:ROM64_INSTR_PT(615) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111111"));
MQQ616:ROM64_INSTR_PT(616) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111111"));
MQQ617:ROM64_INSTR_PT(617) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ618:ROM64_INSTR_PT(618) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ619:ROM64_INSTR_PT(619) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110111"));
MQQ620:ROM64_INSTR_PT(620) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100111"));
MQQ621:ROM64_INSTR_PT(621) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011111"));
MQQ622:ROM64_INSTR_PT(622) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ623:ROM64_INSTR_PT(623) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111111"));
MQQ624:ROM64_INSTR_PT(624) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ625:ROM64_INSTR_PT(625) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ626:ROM64_INSTR_PT(626) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001111"));
MQQ627:ROM64_INSTR_PT(627) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ628:ROM64_INSTR_PT(628) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ629:ROM64_INSTR_PT(629) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ630:ROM64_INSTR_PT(630) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ631:ROM64_INSTR_PT(631) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110011"));
MQQ632:ROM64_INSTR_PT(632) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101011"));
MQQ633:ROM64_INSTR_PT(633) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011011"));
MQQ634:ROM64_INSTR_PT(634) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111011"));
MQQ635:ROM64_INSTR_PT(635) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111011"));
MQQ636:ROM64_INSTR_PT(636) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ637:ROM64_INSTR_PT(637) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ638:ROM64_INSTR_PT(638) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("10011"));
MQQ639:ROM64_INSTR_PT(639) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100111"));
MQQ640:ROM64_INSTR_PT(640) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110111"));
MQQ641:ROM64_INSTR_PT(641) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000111"));
MQQ642:ROM64_INSTR_PT(642) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ643:ROM64_INSTR_PT(643) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ644:ROM64_INSTR_PT(644) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ645:ROM64_INSTR_PT(645) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110111"));
MQQ646:ROM64_INSTR_PT(646) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011111"));
MQQ647:ROM64_INSTR_PT(647) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ648:ROM64_INSTR_PT(648) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ649:ROM64_INSTR_PT(649) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ650:ROM64_INSTR_PT(650) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ651:ROM64_INSTR_PT(651) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("10111"));
MQQ652:ROM64_INSTR_PT(652) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ653:ROM64_INSTR_PT(653) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ654:ROM64_INSTR_PT(654) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000001"));
MQQ655:ROM64_INSTR_PT(655) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110001"));
MQQ656:ROM64_INSTR_PT(656) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110001"));
MQQ657:ROM64_INSTR_PT(657) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101001"));
MQQ658:ROM64_INSTR_PT(658) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001001"));
MQQ659:ROM64_INSTR_PT(659) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011001"));
MQQ660:ROM64_INSTR_PT(660) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101001"));
MQQ661:ROM64_INSTR_PT(661) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000101"));
MQQ662:ROM64_INSTR_PT(662) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000101"));
MQQ663:ROM64_INSTR_PT(663) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100101"));
MQQ664:ROM64_INSTR_PT(664) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110101"));
MQQ665:ROM64_INSTR_PT(665) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001101"));
MQQ666:ROM64_INSTR_PT(666) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011101"));
MQQ667:ROM64_INSTR_PT(667) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011101"));
MQQ668:ROM64_INSTR_PT(668) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000001"));
MQQ669:ROM64_INSTR_PT(669) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010001"));
MQQ670:ROM64_INSTR_PT(670) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110001"));
MQQ671:ROM64_INSTR_PT(671) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001001"));
MQQ672:ROM64_INSTR_PT(672) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0010101"));
MQQ673:ROM64_INSTR_PT(673) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011101"));
MQQ674:ROM64_INSTR_PT(674) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000011"));
MQQ675:ROM64_INSTR_PT(675) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100011"));
MQQ676:ROM64_INSTR_PT(676) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ677:ROM64_INSTR_PT(677) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ678:ROM64_INSTR_PT(678) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101011"));
MQQ679:ROM64_INSTR_PT(679) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011011"));
MQQ680:ROM64_INSTR_PT(680) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011011"));
MQQ681:ROM64_INSTR_PT(681) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ682:ROM64_INSTR_PT(682) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ683:ROM64_INSTR_PT(683) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010011"));
MQQ684:ROM64_INSTR_PT(684) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100111"));
MQQ685:ROM64_INSTR_PT(685) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010111"));
MQQ686:ROM64_INSTR_PT(686) <=
    Eq(( ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0111"));
MQQ687:ROM64_INSTR_PT(687) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001111"));
MQQ688:ROM64_INSTR_PT(688) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101111"));
MQQ689:ROM64_INSTR_PT(689) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011111"));
MQQ690:ROM64_INSTR_PT(690) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ691:ROM64_INSTR_PT(691) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ692:ROM64_INSTR_PT(692) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101111"));
MQQ693:ROM64_INSTR_PT(693) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ694:ROM64_INSTR_PT(694) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000111"));
MQQ695:ROM64_INSTR_PT(695) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110111"));
MQQ696:ROM64_INSTR_PT(696) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("000111"));
MQQ697:ROM64_INSTR_PT(697) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ698:ROM64_INSTR_PT(698) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011111"));
MQQ699:ROM64_INSTR_PT(699) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ700:ROM64_INSTR_PT(700) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011011"));
MQQ701:ROM64_INSTR_PT(701) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ702:ROM64_INSTR_PT(702) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ703:ROM64_INSTR_PT(703) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101111"));
MQQ704:ROM64_INSTR_PT(704) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ705:ROM64_INSTR_PT(705) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ706:ROM64_INSTR_PT(706) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000001"));
MQQ707:ROM64_INSTR_PT(707) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010001"));
MQQ708:ROM64_INSTR_PT(708) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001001"));
MQQ709:ROM64_INSTR_PT(709) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111001"));
MQQ710:ROM64_INSTR_PT(710) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100101"));
MQQ711:ROM64_INSTR_PT(711) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100001"));
MQQ712:ROM64_INSTR_PT(712) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111101"));
MQQ713:ROM64_INSTR_PT(713) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0110111"));
MQQ714:ROM64_INSTR_PT(714) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ715:ROM64_INSTR_PT(715) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ716:ROM64_INSTR_PT(716) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ717:ROM64_INSTR_PT(717) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011111"));
MQQ718:ROM64_INSTR_PT(718) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ719:ROM64_INSTR_PT(719) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100101"));
MQQ720:ROM64_INSTR_PT(720) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ721:ROM64_INSTR_PT(721) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101"));
MQQ722:ROM64_INSTR_PT(722) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100000"));
MQQ723:ROM64_INSTR_PT(723) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100000"));
MQQ724:ROM64_INSTR_PT(724) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("010010000"));
MQQ725:ROM64_INSTR_PT(725) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000110000"));
MQQ726:ROM64_INSTR_PT(726) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ727:ROM64_INSTR_PT(727) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100000"));
MQQ728:ROM64_INSTR_PT(728) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("010001000"));
MQQ729:ROM64_INSTR_PT(729) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11011000"));
MQQ730:ROM64_INSTR_PT(730) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111000"));
MQQ731:ROM64_INSTR_PT(731) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0111000"));
MQQ732:ROM64_INSTR_PT(732) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110000"));
MQQ733:ROM64_INSTR_PT(733) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00000100"));
MQQ734:ROM64_INSTR_PT(734) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000100"));
MQQ735:ROM64_INSTR_PT(735) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100100"));
MQQ736:ROM64_INSTR_PT(736) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1100100"));
MQQ737:ROM64_INSTR_PT(737) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100100"));
MQQ738:ROM64_INSTR_PT(738) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("010010100"));
MQQ739:ROM64_INSTR_PT(739) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ740:ROM64_INSTR_PT(740) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ741:ROM64_INSTR_PT(741) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("10011100"));
MQQ742:ROM64_INSTR_PT(742) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101100"));
MQQ743:ROM64_INSTR_PT(743) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0111100"));
MQQ744:ROM64_INSTR_PT(744) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100100"));
MQQ745:ROM64_INSTR_PT(745) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100000"));
MQQ746:ROM64_INSTR_PT(746) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1100000"));
MQQ747:ROM64_INSTR_PT(747) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00000100"));
MQQ748:ROM64_INSTR_PT(748) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0101100"));
MQQ749:ROM64_INSTR_PT(749) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011100"));
MQQ750:ROM64_INSTR_PT(750) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ751:ROM64_INSTR_PT(751) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11100"));
MQQ752:ROM64_INSTR_PT(752) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000"));
MQQ753:ROM64_INSTR_PT(753) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100010"));
MQQ754:ROM64_INSTR_PT(754) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00010010"));
MQQ755:ROM64_INSTR_PT(755) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00000010"));
MQQ756:ROM64_INSTR_PT(756) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11001010"));
MQQ757:ROM64_INSTR_PT(757) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111010"));
MQQ758:ROM64_INSTR_PT(758) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1111010"));
MQQ759:ROM64_INSTR_PT(759) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101010"));
MQQ760:ROM64_INSTR_PT(760) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1000110"));
MQQ761:ROM64_INSTR_PT(761) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("110100110"));
MQQ762:ROM64_INSTR_PT(762) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0010110"));
MQQ763:ROM64_INSTR_PT(763) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("010110"));
MQQ764:ROM64_INSTR_PT(764) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0001110"));
MQQ765:ROM64_INSTR_PT(765) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011110"));
MQQ766:ROM64_INSTR_PT(766) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("10011110"));
MQQ767:ROM64_INSTR_PT(767) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ768:ROM64_INSTR_PT(768) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("0110"));
MQQ769:ROM64_INSTR_PT(769) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011110"));
MQQ770:ROM64_INSTR_PT(770) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ771:ROM64_INSTR_PT(771) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("010110"));
MQQ772:ROM64_INSTR_PT(772) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("10000"));
MQQ773:ROM64_INSTR_PT(773) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ774:ROM64_INSTR_PT(774) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011100"));
MQQ775:ROM64_INSTR_PT(775) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("00100"));
MQQ776:ROM64_INSTR_PT(776) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100010"));
MQQ777:ROM64_INSTR_PT(777) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11010010"));
MQQ778:ROM64_INSTR_PT(778) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101010"));
MQQ779:ROM64_INSTR_PT(779) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01110"));
MQQ780:ROM64_INSTR_PT(780) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01110"));
MQQ781:ROM64_INSTR_PT(781) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01000001"));
MQQ782:ROM64_INSTR_PT(782) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("110100001"));
MQQ783:ROM64_INSTR_PT(783) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01010001"));
MQQ784:ROM64_INSTR_PT(784) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11010001"));
MQQ785:ROM64_INSTR_PT(785) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1010001"));
MQQ786:ROM64_INSTR_PT(786) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000001"));
MQQ787:ROM64_INSTR_PT(787) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("010001"));
MQQ788:ROM64_INSTR_PT(788) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0001001"));
MQQ789:ROM64_INSTR_PT(789) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("001001"));
MQQ790:ROM64_INSTR_PT(790) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011001"));
MQQ791:ROM64_INSTR_PT(791) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111001"));
MQQ792:ROM64_INSTR_PT(792) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011001"));
MQQ793:ROM64_INSTR_PT(793) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111001"));
MQQ794:ROM64_INSTR_PT(794) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00100101"));
MQQ795:ROM64_INSTR_PT(795) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00010101"));
MQQ796:ROM64_INSTR_PT(796) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011101"));
MQQ797:ROM64_INSTR_PT(797) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("10011101"));
MQQ798:ROM64_INSTR_PT(798) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110101"));
MQQ799:ROM64_INSTR_PT(799) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("10101"));
MQQ800:ROM64_INSTR_PT(800) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11101"));
MQQ801:ROM64_INSTR_PT(801) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000101"));
MQQ802:ROM64_INSTR_PT(802) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000101"));
MQQ803:ROM64_INSTR_PT(803) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11101"));
MQQ804:ROM64_INSTR_PT(804) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000100011"));
MQQ805:ROM64_INSTR_PT(805) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01110011"));
MQQ806:ROM64_INSTR_PT(806) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00000011"));
MQQ807:ROM64_INSTR_PT(807) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000011"));
MQQ808:ROM64_INSTR_PT(808) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000011"));
MQQ809:ROM64_INSTR_PT(809) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1010011"));
MQQ810:ROM64_INSTR_PT(810) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("010011"));
MQQ811:ROM64_INSTR_PT(811) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01101011"));
MQQ812:ROM64_INSTR_PT(812) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00001011"));
MQQ813:ROM64_INSTR_PT(813) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ814:ROM64_INSTR_PT(814) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101011"));
MQQ815:ROM64_INSTR_PT(815) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ816:ROM64_INSTR_PT(816) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100111"));
MQQ817:ROM64_INSTR_PT(817) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00010111"));
MQQ818:ROM64_INSTR_PT(818) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ819:ROM64_INSTR_PT(819) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1110111"));
MQQ820:ROM64_INSTR_PT(820) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11010111"));
MQQ821:ROM64_INSTR_PT(821) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000101111"));
MQQ822:ROM64_INSTR_PT(822) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01101111"));
MQQ823:ROM64_INSTR_PT(823) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ824:ROM64_INSTR_PT(824) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ825:ROM64_INSTR_PT(825) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ826:ROM64_INSTR_PT(826) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ827:ROM64_INSTR_PT(827) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101011"));
MQQ828:ROM64_INSTR_PT(828) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0110111"));
MQQ829:ROM64_INSTR_PT(829) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ830:ROM64_INSTR_PT(830) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ831:ROM64_INSTR_PT(831) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("0111"));
MQQ832:ROM64_INSTR_PT(832) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ833:ROM64_INSTR_PT(833) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ834:ROM64_INSTR_PT(834) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110001"));
MQQ835:ROM64_INSTR_PT(835) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1001101"));
MQQ836:ROM64_INSTR_PT(836) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101101"));
MQQ837:ROM64_INSTR_PT(837) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101011"));
MQQ838:ROM64_INSTR_PT(838) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1111011"));
MQQ839:ROM64_INSTR_PT(839) <=
    Eq(( ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("011"));
MQQ840:ROM64_INSTR_PT(840) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000111"));
MQQ841:ROM64_INSTR_PT(841) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ842:ROM64_INSTR_PT(842) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101111"));
MQQ843:ROM64_INSTR_PT(843) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01111"));
MQQ844:ROM64_INSTR_PT(844) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ845:ROM64_INSTR_PT(845) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ846:ROM64_INSTR_PT(846) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011111"));
MQQ847:ROM64_INSTR_PT(847) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("000101"));
MQQ848:ROM64_INSTR_PT(848) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01101"));
MQQ849:ROM64_INSTR_PT(849) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ850:ROM64_INSTR_PT(850) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("1111"));
MQQ851:ROM64_INSTR_PT(851) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01001"));
MQQ852:ROM64_INSTR_PT(852) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1001000"));
MQQ853:ROM64_INSTR_PT(853) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("110000"));
MQQ854:ROM64_INSTR_PT(854) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("00011100"));
MQQ855:ROM64_INSTR_PT(855) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("00000010"));
MQQ856:ROM64_INSTR_PT(856) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0100010"));
MQQ857:ROM64_INSTR_PT(857) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0000010"));
MQQ858:ROM64_INSTR_PT(858) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("101110"));
MQQ859:ROM64_INSTR_PT(859) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1101110"));
MQQ860:ROM64_INSTR_PT(860) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("000110"));
MQQ861:ROM64_INSTR_PT(861) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1001100"));
MQQ862:ROM64_INSTR_PT(862) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("1110"));
MQQ863:ROM64_INSTR_PT(863) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("010"));
MQQ864:ROM64_INSTR_PT(864) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0100101"));
MQQ865:ROM64_INSTR_PT(865) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1100101"));
MQQ866:ROM64_INSTR_PT(866) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1001101"));
MQQ867:ROM64_INSTR_PT(867) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1101101"));
MQQ868:ROM64_INSTR_PT(868) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("01011"));
MQQ869:ROM64_INSTR_PT(869) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ870:ROM64_INSTR_PT(870) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0011111"));
MQQ871:ROM64_INSTR_PT(871) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("100111"));
MQQ872:ROM64_INSTR_PT(872) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ873:ROM64_INSTR_PT(873) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ874:ROM64_INSTR_PT(874) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ875:ROM64_INSTR_PT(875) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("01111"));
MQQ876:ROM64_INSTR_PT(876) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("101"));
MQQ877:ROM64_INSTR_PT(877) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("010001"));
MQQ878:ROM64_INSTR_PT(878) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("01111"));
MQQ879:ROM64_INSTR_PT(879) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("111"));
MQQ880:ROM64_INSTR_PT(880) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) ) , STD_ULOGIC_VECTOR'("01110"));
MQQ881:ROM64_INSTR_PT(881) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(6)
     ) , STD_ULOGIC_VECTOR'("00"));
MQQ882:ROM64_INSTR_PT(882) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) ) , STD_ULOGIC_VECTOR'("111"));
MQQ883:ROM64_INSTR_PT(883) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ884:ROM64_INSTR_PT(884) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5)
     ) , STD_ULOGIC_VECTOR'("00"));
MQQ885:ROM64_INSTR_PT(885) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) ) , STD_ULOGIC_VECTOR'("111"));
MQQ886:ROM64_INSTR_PT(886) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) ) , STD_ULOGIC_VECTOR'("111"));
MQQ887:ROM64_INSTR_PT(887) <=
    Eq(( ROM_ADDR_L2(2) ) , STD_ULOGIC'('1'));
MQQ888:ROM64_INSTR_PT(888) <=
    Eq(( ROM_ADDR_L2(1) ) , STD_ULOGIC'('1'));
MQQ889:ROM64_INSTR_PT(889) <=
    Eq(( ROM_ADDR_L2(0) ) , STD_ULOGIC'('0'));
MQQ890:ROM64_INSTR_PT(890) <=
    '1';
MQQ891:TEMPLATE(0) <= 
    (ROM64_INSTR_PT(29) OR ROM64_INSTR_PT(35)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(65)
     OR ROM64_INSTR_PT(74) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(112) OR ROM64_INSTR_PT(119)
     OR ROM64_INSTR_PT(129) OR ROM64_INSTR_PT(134)
     OR ROM64_INSTR_PT(143) OR ROM64_INSTR_PT(158)
     OR ROM64_INSTR_PT(160) OR ROM64_INSTR_PT(176)
     OR ROM64_INSTR_PT(177) OR ROM64_INSTR_PT(179)
     OR ROM64_INSTR_PT(183) OR ROM64_INSTR_PT(221)
     OR ROM64_INSTR_PT(225) OR ROM64_INSTR_PT(233)
     OR ROM64_INSTR_PT(237) OR ROM64_INSTR_PT(242)
     OR ROM64_INSTR_PT(259) OR ROM64_INSTR_PT(294)
     OR ROM64_INSTR_PT(296) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(339) OR ROM64_INSTR_PT(350)
     OR ROM64_INSTR_PT(354) OR ROM64_INSTR_PT(355)
     OR ROM64_INSTR_PT(358) OR ROM64_INSTR_PT(359)
     OR ROM64_INSTR_PT(362) OR ROM64_INSTR_PT(367)
     OR ROM64_INSTR_PT(368) OR ROM64_INSTR_PT(378)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(389)
     OR ROM64_INSTR_PT(392) OR ROM64_INSTR_PT(402)
     OR ROM64_INSTR_PT(428) OR ROM64_INSTR_PT(435)
     OR ROM64_INSTR_PT(470) OR ROM64_INSTR_PT(477)
     OR ROM64_INSTR_PT(527) OR ROM64_INSTR_PT(557)
     OR ROM64_INSTR_PT(564) OR ROM64_INSTR_PT(572)
     OR ROM64_INSTR_PT(590) OR ROM64_INSTR_PT(602)
     OR ROM64_INSTR_PT(610) OR ROM64_INSTR_PT(619)
     OR ROM64_INSTR_PT(653) OR ROM64_INSTR_PT(657)
     OR ROM64_INSTR_PT(664) OR ROM64_INSTR_PT(694)
     OR ROM64_INSTR_PT(695) OR ROM64_INSTR_PT(702)
     OR ROM64_INSTR_PT(716) OR ROM64_INSTR_PT(719)
     OR ROM64_INSTR_PT(720) OR ROM64_INSTR_PT(721)
     OR ROM64_INSTR_PT(736) OR ROM64_INSTR_PT(770)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(832)
     OR ROM64_INSTR_PT(834) OR ROM64_INSTR_PT(858)
     OR ROM64_INSTR_PT(873));
MQQ892:TEMPLATE(1) <= 
    (ROM64_INSTR_PT(2) OR ROM64_INSTR_PT(4)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(8)
     OR ROM64_INSTR_PT(9) OR ROM64_INSTR_PT(10)
     OR ROM64_INSTR_PT(11) OR ROM64_INSTR_PT(14)
     OR ROM64_INSTR_PT(15) OR ROM64_INSTR_PT(17)
     OR ROM64_INSTR_PT(18) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(25)
     OR ROM64_INSTR_PT(34) OR ROM64_INSTR_PT(36)
     OR ROM64_INSTR_PT(38) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(43)
     OR ROM64_INSTR_PT(49) OR ROM64_INSTR_PT(51)
     OR ROM64_INSTR_PT(52) OR ROM64_INSTR_PT(53)
     OR ROM64_INSTR_PT(55) OR ROM64_INSTR_PT(56)
     OR ROM64_INSTR_PT(61) OR ROM64_INSTR_PT(64)
     OR ROM64_INSTR_PT(68) OR ROM64_INSTR_PT(69)
     OR ROM64_INSTR_PT(70) OR ROM64_INSTR_PT(71)
     OR ROM64_INSTR_PT(73) OR ROM64_INSTR_PT(75)
     OR ROM64_INSTR_PT(77) OR ROM64_INSTR_PT(78)
     OR ROM64_INSTR_PT(82) OR ROM64_INSTR_PT(83)
     OR ROM64_INSTR_PT(86) OR ROM64_INSTR_PT(89)
     OR ROM64_INSTR_PT(90) OR ROM64_INSTR_PT(92)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(95)
     OR ROM64_INSTR_PT(96) OR ROM64_INSTR_PT(97)
     OR ROM64_INSTR_PT(99) OR ROM64_INSTR_PT(100)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(102)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(105)
     OR ROM64_INSTR_PT(106) OR ROM64_INSTR_PT(108)
     OR ROM64_INSTR_PT(109) OR ROM64_INSTR_PT(110)
     OR ROM64_INSTR_PT(113) OR ROM64_INSTR_PT(116)
     OR ROM64_INSTR_PT(117) OR ROM64_INSTR_PT(118)
     OR ROM64_INSTR_PT(124) OR ROM64_INSTR_PT(127)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(144)
     OR ROM64_INSTR_PT(145) OR ROM64_INSTR_PT(148)
     OR ROM64_INSTR_PT(153) OR ROM64_INSTR_PT(161)
     OR ROM64_INSTR_PT(162) OR ROM64_INSTR_PT(164)
     OR ROM64_INSTR_PT(169) OR ROM64_INSTR_PT(170)
     OR ROM64_INSTR_PT(171) OR ROM64_INSTR_PT(172)
     OR ROM64_INSTR_PT(173) OR ROM64_INSTR_PT(175)
     OR ROM64_INSTR_PT(180) OR ROM64_INSTR_PT(184)
     OR ROM64_INSTR_PT(185) OR ROM64_INSTR_PT(186)
     OR ROM64_INSTR_PT(188) OR ROM64_INSTR_PT(193)
     OR ROM64_INSTR_PT(195) OR ROM64_INSTR_PT(196)
     OR ROM64_INSTR_PT(199) OR ROM64_INSTR_PT(201)
     OR ROM64_INSTR_PT(202) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(205) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(208) OR ROM64_INSTR_PT(214)
     OR ROM64_INSTR_PT(215) OR ROM64_INSTR_PT(216)
     OR ROM64_INSTR_PT(217) OR ROM64_INSTR_PT(218)
     OR ROM64_INSTR_PT(222) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(226) OR ROM64_INSTR_PT(229)
     OR ROM64_INSTR_PT(230) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(241) OR ROM64_INSTR_PT(243)
     OR ROM64_INSTR_PT(244) OR ROM64_INSTR_PT(252)
     OR ROM64_INSTR_PT(254) OR ROM64_INSTR_PT(257)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(263)
     OR ROM64_INSTR_PT(264) OR ROM64_INSTR_PT(265)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(269)
     OR ROM64_INSTR_PT(270) OR ROM64_INSTR_PT(271)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(275)
     OR ROM64_INSTR_PT(276) OR ROM64_INSTR_PT(277)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(282)
     OR ROM64_INSTR_PT(284) OR ROM64_INSTR_PT(285)
     OR ROM64_INSTR_PT(286) OR ROM64_INSTR_PT(287)
     OR ROM64_INSTR_PT(292) OR ROM64_INSTR_PT(293)
     OR ROM64_INSTR_PT(297) OR ROM64_INSTR_PT(298)
     OR ROM64_INSTR_PT(299) OR ROM64_INSTR_PT(302)
     OR ROM64_INSTR_PT(305) OR ROM64_INSTR_PT(308)
     OR ROM64_INSTR_PT(315) OR ROM64_INSTR_PT(322)
     OR ROM64_INSTR_PT(325) OR ROM64_INSTR_PT(331)
     OR ROM64_INSTR_PT(333) OR ROM64_INSTR_PT(345)
     OR ROM64_INSTR_PT(349) OR ROM64_INSTR_PT(351)
     OR ROM64_INSTR_PT(357) OR ROM64_INSTR_PT(364)
     OR ROM64_INSTR_PT(365) OR ROM64_INSTR_PT(366)
     OR ROM64_INSTR_PT(369) OR ROM64_INSTR_PT(371)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(375)
     OR ROM64_INSTR_PT(377) OR ROM64_INSTR_PT(379)
     OR ROM64_INSTR_PT(381) OR ROM64_INSTR_PT(383)
     OR ROM64_INSTR_PT(385) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(391) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(403) OR ROM64_INSTR_PT(404)
     OR ROM64_INSTR_PT(405) OR ROM64_INSTR_PT(408)
     OR ROM64_INSTR_PT(409) OR ROM64_INSTR_PT(410)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(419) OR ROM64_INSTR_PT(420)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(424)
     OR ROM64_INSTR_PT(425) OR ROM64_INSTR_PT(426)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(429)
     OR ROM64_INSTR_PT(430) OR ROM64_INSTR_PT(432)
     OR ROM64_INSTR_PT(433) OR ROM64_INSTR_PT(434)
     OR ROM64_INSTR_PT(437) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(439) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(443) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(451)
     OR ROM64_INSTR_PT(453) OR ROM64_INSTR_PT(454)
     OR ROM64_INSTR_PT(455) OR ROM64_INSTR_PT(456)
     OR ROM64_INSTR_PT(457) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(460) OR ROM64_INSTR_PT(463)
     OR ROM64_INSTR_PT(466) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(478) OR ROM64_INSTR_PT(480)
     OR ROM64_INSTR_PT(481) OR ROM64_INSTR_PT(482)
     OR ROM64_INSTR_PT(483) OR ROM64_INSTR_PT(484)
     OR ROM64_INSTR_PT(485) OR ROM64_INSTR_PT(490)
     OR ROM64_INSTR_PT(493) OR ROM64_INSTR_PT(495)
     OR ROM64_INSTR_PT(497) OR ROM64_INSTR_PT(498)
     OR ROM64_INSTR_PT(499) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(505)
     OR ROM64_INSTR_PT(506) OR ROM64_INSTR_PT(508)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(510)
     OR ROM64_INSTR_PT(511) OR ROM64_INSTR_PT(512)
     OR ROM64_INSTR_PT(514) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(521) OR ROM64_INSTR_PT(522)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(525)
     OR ROM64_INSTR_PT(530) OR ROM64_INSTR_PT(531)
     OR ROM64_INSTR_PT(532) OR ROM64_INSTR_PT(534)
     OR ROM64_INSTR_PT(535) OR ROM64_INSTR_PT(536)
     OR ROM64_INSTR_PT(537) OR ROM64_INSTR_PT(539)
     OR ROM64_INSTR_PT(540) OR ROM64_INSTR_PT(542)
     OR ROM64_INSTR_PT(544) OR ROM64_INSTR_PT(545)
     OR ROM64_INSTR_PT(546) OR ROM64_INSTR_PT(548)
     OR ROM64_INSTR_PT(549) OR ROM64_INSTR_PT(552)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(555) OR ROM64_INSTR_PT(558)
     OR ROM64_INSTR_PT(559) OR ROM64_INSTR_PT(563)
     OR ROM64_INSTR_PT(566) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(569) OR ROM64_INSTR_PT(570)
     OR ROM64_INSTR_PT(571) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(577)
     OR ROM64_INSTR_PT(579) OR ROM64_INSTR_PT(580)
     OR ROM64_INSTR_PT(581) OR ROM64_INSTR_PT(582)
     OR ROM64_INSTR_PT(583) OR ROM64_INSTR_PT(584)
     OR ROM64_INSTR_PT(586) OR ROM64_INSTR_PT(588)
     OR ROM64_INSTR_PT(589) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(592) OR ROM64_INSTR_PT(593)
     OR ROM64_INSTR_PT(595) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(598) OR ROM64_INSTR_PT(599)
     OR ROM64_INSTR_PT(600) OR ROM64_INSTR_PT(603)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(606)
     OR ROM64_INSTR_PT(607) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(611) OR ROM64_INSTR_PT(612)
     OR ROM64_INSTR_PT(613) OR ROM64_INSTR_PT(614)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(616)
     OR ROM64_INSTR_PT(617) OR ROM64_INSTR_PT(618)
     OR ROM64_INSTR_PT(623) OR ROM64_INSTR_PT(626)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(629) OR ROM64_INSTR_PT(633)
     OR ROM64_INSTR_PT(637) OR ROM64_INSTR_PT(639)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(643)
     OR ROM64_INSTR_PT(644) OR ROM64_INSTR_PT(646)
     OR ROM64_INSTR_PT(655) OR ROM64_INSTR_PT(660)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(666)
     OR ROM64_INSTR_PT(678) OR ROM64_INSTR_PT(679)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(682)
     OR ROM64_INSTR_PT(687) OR ROM64_INSTR_PT(703)
     OR ROM64_INSTR_PT(713) OR ROM64_INSTR_PT(717)
     OR ROM64_INSTR_PT(722) OR ROM64_INSTR_PT(731)
     OR ROM64_INSTR_PT(741) OR ROM64_INSTR_PT(744)
     OR ROM64_INSTR_PT(753) OR ROM64_INSTR_PT(761)
     OR ROM64_INSTR_PT(769) OR ROM64_INSTR_PT(776)
     OR ROM64_INSTR_PT(791) OR ROM64_INSTR_PT(801)
     OR ROM64_INSTR_PT(808) OR ROM64_INSTR_PT(811)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(822)
     OR ROM64_INSTR_PT(824) OR ROM64_INSTR_PT(846)
     OR ROM64_INSTR_PT(849) OR ROM64_INSTR_PT(852)
     OR ROM64_INSTR_PT(854) OR ROM64_INSTR_PT(855)
     OR ROM64_INSTR_PT(856) OR ROM64_INSTR_PT(864)
     OR ROM64_INSTR_PT(869) OR ROM64_INSTR_PT(870)
     OR ROM64_INSTR_PT(872) OR ROM64_INSTR_PT(886)
    );
MQQ893:TEMPLATE(2) <= 
    (ROM64_INSTR_PT(2) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(10)
     OR ROM64_INSTR_PT(14) OR ROM64_INSTR_PT(15)
     OR ROM64_INSTR_PT(18) OR ROM64_INSTR_PT(20)
     OR ROM64_INSTR_PT(25) OR ROM64_INSTR_PT(28)
     OR ROM64_INSTR_PT(33) OR ROM64_INSTR_PT(36)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(43)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(56)
     OR ROM64_INSTR_PT(60) OR ROM64_INSTR_PT(66)
     OR ROM64_INSTR_PT(69) OR ROM64_INSTR_PT(73)
     OR ROM64_INSTR_PT(77) OR ROM64_INSTR_PT(78)
     OR ROM64_INSTR_PT(79) OR ROM64_INSTR_PT(82)
     OR ROM64_INSTR_PT(89) OR ROM64_INSTR_PT(92)
     OR ROM64_INSTR_PT(95) OR ROM64_INSTR_PT(96)
     OR ROM64_INSTR_PT(97) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(104)
     OR ROM64_INSTR_PT(106) OR ROM64_INSTR_PT(108)
     OR ROM64_INSTR_PT(109) OR ROM64_INSTR_PT(110)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(124)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(142)
     OR ROM64_INSTR_PT(145) OR ROM64_INSTR_PT(146)
     OR ROM64_INSTR_PT(147) OR ROM64_INSTR_PT(150)
     OR ROM64_INSTR_PT(151) OR ROM64_INSTR_PT(153)
     OR ROM64_INSTR_PT(161) OR ROM64_INSTR_PT(166)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(172)
     OR ROM64_INSTR_PT(173) OR ROM64_INSTR_PT(174)
     OR ROM64_INSTR_PT(175) OR ROM64_INSTR_PT(184)
     OR ROM64_INSTR_PT(187) OR ROM64_INSTR_PT(188)
     OR ROM64_INSTR_PT(190) OR ROM64_INSTR_PT(191)
     OR ROM64_INSTR_PT(193) OR ROM64_INSTR_PT(195)
     OR ROM64_INSTR_PT(202) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(205) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(207) OR ROM64_INSTR_PT(208)
     OR ROM64_INSTR_PT(209) OR ROM64_INSTR_PT(216)
     OR ROM64_INSTR_PT(219) OR ROM64_INSTR_PT(228)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(231) OR ROM64_INSTR_PT(240)
     OR ROM64_INSTR_PT(243) OR ROM64_INSTR_PT(247)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(254)
     OR ROM64_INSTR_PT(257) OR ROM64_INSTR_PT(258)
     OR ROM64_INSTR_PT(260) OR ROM64_INSTR_PT(261)
     OR ROM64_INSTR_PT(265) OR ROM64_INSTR_PT(269)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(277)
     OR ROM64_INSTR_PT(281) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(288) OR ROM64_INSTR_PT(292)
     OR ROM64_INSTR_PT(295) OR ROM64_INSTR_PT(304)
     OR ROM64_INSTR_PT(307) OR ROM64_INSTR_PT(309)
     OR ROM64_INSTR_PT(313) OR ROM64_INSTR_PT(324)
     OR ROM64_INSTR_PT(325) OR ROM64_INSTR_PT(327)
     OR ROM64_INSTR_PT(332) OR ROM64_INSTR_PT(333)
     OR ROM64_INSTR_PT(334) OR ROM64_INSTR_PT(340)
     OR ROM64_INSTR_PT(341) OR ROM64_INSTR_PT(342)
     OR ROM64_INSTR_PT(345) OR ROM64_INSTR_PT(351)
     OR ROM64_INSTR_PT(352) OR ROM64_INSTR_PT(357)
     OR ROM64_INSTR_PT(361) OR ROM64_INSTR_PT(365)
     OR ROM64_INSTR_PT(366) OR ROM64_INSTR_PT(369)
     OR ROM64_INSTR_PT(371) OR ROM64_INSTR_PT(372)
     OR ROM64_INSTR_PT(374) OR ROM64_INSTR_PT(377)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(388) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(396)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(403)
     OR ROM64_INSTR_PT(405) OR ROM64_INSTR_PT(406)
     OR ROM64_INSTR_PT(408) OR ROM64_INSTR_PT(409)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(419) OR ROM64_INSTR_PT(420)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(425)
     OR ROM64_INSTR_PT(426) OR ROM64_INSTR_PT(429)
     OR ROM64_INSTR_PT(430) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(439) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(443) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(448)
     OR ROM64_INSTR_PT(451) OR ROM64_INSTR_PT(453)
     OR ROM64_INSTR_PT(454) OR ROM64_INSTR_PT(455)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(460) OR ROM64_INSTR_PT(463)
     OR ROM64_INSTR_PT(464) OR ROM64_INSTR_PT(466)
     OR ROM64_INSTR_PT(467) OR ROM64_INSTR_PT(468)
     OR ROM64_INSTR_PT(471) OR ROM64_INSTR_PT(472)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(474)
     OR ROM64_INSTR_PT(475) OR ROM64_INSTR_PT(483)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(491)
     OR ROM64_INSTR_PT(497) OR ROM64_INSTR_PT(498)
     OR ROM64_INSTR_PT(499) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(506) OR ROM64_INSTR_PT(508)
     OR ROM64_INSTR_PT(510) OR ROM64_INSTR_PT(514)
     OR ROM64_INSTR_PT(516) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(532) OR ROM64_INSTR_PT(538)
     OR ROM64_INSTR_PT(542) OR ROM64_INSTR_PT(546)
     OR ROM64_INSTR_PT(549) OR ROM64_INSTR_PT(551)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(559) OR ROM64_INSTR_PT(562)
     OR ROM64_INSTR_PT(566) OR ROM64_INSTR_PT(570)
     OR ROM64_INSTR_PT(571) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(581)
     OR ROM64_INSTR_PT(586) OR ROM64_INSTR_PT(589)
     OR ROM64_INSTR_PT(593) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(598)
     OR ROM64_INSTR_PT(601) OR ROM64_INSTR_PT(603)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(606)
     OR ROM64_INSTR_PT(611) OR ROM64_INSTR_PT(612)
     OR ROM64_INSTR_PT(613) OR ROM64_INSTR_PT(614)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(616)
     OR ROM64_INSTR_PT(617) OR ROM64_INSTR_PT(620)
     OR ROM64_INSTR_PT(626) OR ROM64_INSTR_PT(627)
     OR ROM64_INSTR_PT(628) OR ROM64_INSTR_PT(632)
     OR ROM64_INSTR_PT(635) OR ROM64_INSTR_PT(654)
     OR ROM64_INSTR_PT(659) OR ROM64_INSTR_PT(660)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(668)
     OR ROM64_INSTR_PT(675) OR ROM64_INSTR_PT(679)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(682)
     OR ROM64_INSTR_PT(687) OR ROM64_INSTR_PT(691)
     OR ROM64_INSTR_PT(703) OR ROM64_INSTR_PT(709)
     OR ROM64_INSTR_PT(711) OR ROM64_INSTR_PT(713)
     OR ROM64_INSTR_PT(717) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(728)
     OR ROM64_INSTR_PT(733) OR ROM64_INSTR_PT(735)
     OR ROM64_INSTR_PT(738) OR ROM64_INSTR_PT(741)
     OR ROM64_INSTR_PT(759) OR ROM64_INSTR_PT(766)
     OR ROM64_INSTR_PT(781) OR ROM64_INSTR_PT(791)
     OR ROM64_INSTR_PT(794) OR ROM64_INSTR_PT(797)
     OR ROM64_INSTR_PT(801) OR ROM64_INSTR_PT(808)
     OR ROM64_INSTR_PT(809) OR ROM64_INSTR_PT(811)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(822)
     OR ROM64_INSTR_PT(824) OR ROM64_INSTR_PT(846)
     OR ROM64_INSTR_PT(849) OR ROM64_INSTR_PT(852)
     OR ROM64_INSTR_PT(854) OR ROM64_INSTR_PT(855)
     OR ROM64_INSTR_PT(869) OR ROM64_INSTR_PT(872)
     OR ROM64_INSTR_PT(883) OR ROM64_INSTR_PT(886)
    );
MQQ894:TEMPLATE(3) <= 
    (ROM64_INSTR_PT(2) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(9)
     OR ROM64_INSTR_PT(10) OR ROM64_INSTR_PT(11)
     OR ROM64_INSTR_PT(14) OR ROM64_INSTR_PT(15)
     OR ROM64_INSTR_PT(17) OR ROM64_INSTR_PT(18)
     OR ROM64_INSTR_PT(20) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(25)
     OR ROM64_INSTR_PT(28) OR ROM64_INSTR_PT(29)
     OR ROM64_INSTR_PT(33) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(35) OR ROM64_INSTR_PT(36)
     OR ROM64_INSTR_PT(38) OR ROM64_INSTR_PT(39)
     OR ROM64_INSTR_PT(41) OR ROM64_INSTR_PT(42)
     OR ROM64_INSTR_PT(43) OR ROM64_INSTR_PT(45)
     OR ROM64_INSTR_PT(49) OR ROM64_INSTR_PT(52)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(56)
     OR ROM64_INSTR_PT(60) OR ROM64_INSTR_PT(61)
     OR ROM64_INSTR_PT(64) OR ROM64_INSTR_PT(66)
     OR ROM64_INSTR_PT(69) OR ROM64_INSTR_PT(70)
     OR ROM64_INSTR_PT(71) OR ROM64_INSTR_PT(73)
     OR ROM64_INSTR_PT(75) OR ROM64_INSTR_PT(76)
     OR ROM64_INSTR_PT(77) OR ROM64_INSTR_PT(78)
     OR ROM64_INSTR_PT(80) OR ROM64_INSTR_PT(82)
     OR ROM64_INSTR_PT(83) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(86) OR ROM64_INSTR_PT(89)
     OR ROM64_INSTR_PT(90) OR ROM64_INSTR_PT(92)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(95)
     OR ROM64_INSTR_PT(96) OR ROM64_INSTR_PT(97)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(99)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(102)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(106)
     OR ROM64_INSTR_PT(108) OR ROM64_INSTR_PT(109)
     OR ROM64_INSTR_PT(110) OR ROM64_INSTR_PT(113)
     OR ROM64_INSTR_PT(114) OR ROM64_INSTR_PT(115)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(124)
     OR ROM64_INSTR_PT(127) OR ROM64_INSTR_PT(133)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(140)
     OR ROM64_INSTR_PT(142) OR ROM64_INSTR_PT(144)
     OR ROM64_INSTR_PT(145) OR ROM64_INSTR_PT(146)
     OR ROM64_INSTR_PT(147) OR ROM64_INSTR_PT(148)
     OR ROM64_INSTR_PT(150) OR ROM64_INSTR_PT(151)
     OR ROM64_INSTR_PT(153) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(160) OR ROM64_INSTR_PT(161)
     OR ROM64_INSTR_PT(164) OR ROM64_INSTR_PT(166)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(169)
     OR ROM64_INSTR_PT(171) OR ROM64_INSTR_PT(172)
     OR ROM64_INSTR_PT(173) OR ROM64_INSTR_PT(174)
     OR ROM64_INSTR_PT(175) OR ROM64_INSTR_PT(177)
     OR ROM64_INSTR_PT(179) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(181) OR ROM64_INSTR_PT(182)
     OR ROM64_INSTR_PT(183) OR ROM64_INSTR_PT(184)
     OR ROM64_INSTR_PT(186) OR ROM64_INSTR_PT(187)
     OR ROM64_INSTR_PT(188) OR ROM64_INSTR_PT(191)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(199)
     OR ROM64_INSTR_PT(201) OR ROM64_INSTR_PT(202)
     OR ROM64_INSTR_PT(203) OR ROM64_INSTR_PT(205)
     OR ROM64_INSTR_PT(206) OR ROM64_INSTR_PT(207)
     OR ROM64_INSTR_PT(208) OR ROM64_INSTR_PT(209)
     OR ROM64_INSTR_PT(211) OR ROM64_INSTR_PT(215)
     OR ROM64_INSTR_PT(216) OR ROM64_INSTR_PT(217)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(219)
     OR ROM64_INSTR_PT(221) OR ROM64_INSTR_PT(222)
     OR ROM64_INSTR_PT(223) OR ROM64_INSTR_PT(225)
     OR ROM64_INSTR_PT(226) OR ROM64_INSTR_PT(228)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(231) OR ROM64_INSTR_PT(233)
     OR ROM64_INSTR_PT(238) OR ROM64_INSTR_PT(240)
     OR ROM64_INSTR_PT(242) OR ROM64_INSTR_PT(243)
     OR ROM64_INSTR_PT(245) OR ROM64_INSTR_PT(247)
     OR ROM64_INSTR_PT(249) OR ROM64_INSTR_PT(252)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(254)
     OR ROM64_INSTR_PT(257) OR ROM64_INSTR_PT(258)
     OR ROM64_INSTR_PT(259) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(265) OR ROM64_INSTR_PT(268)
     OR ROM64_INSTR_PT(269) OR ROM64_INSTR_PT(270)
     OR ROM64_INSTR_PT(271) OR ROM64_INSTR_PT(272)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(274)
     OR ROM64_INSTR_PT(275) OR ROM64_INSTR_PT(277)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(281)
     OR ROM64_INSTR_PT(282) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(287) OR ROM64_INSTR_PT(288)
     OR ROM64_INSTR_PT(290) OR ROM64_INSTR_PT(293)
     OR ROM64_INSTR_PT(294) OR ROM64_INSTR_PT(295)
     OR ROM64_INSTR_PT(298) OR ROM64_INSTR_PT(299)
     OR ROM64_INSTR_PT(302) OR ROM64_INSTR_PT(304)
     OR ROM64_INSTR_PT(305) OR ROM64_INSTR_PT(307)
     OR ROM64_INSTR_PT(309) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(313) OR ROM64_INSTR_PT(315)
     OR ROM64_INSTR_PT(319) OR ROM64_INSTR_PT(324)
     OR ROM64_INSTR_PT(325) OR ROM64_INSTR_PT(327)
     OR ROM64_INSTR_PT(331) OR ROM64_INSTR_PT(332)
     OR ROM64_INSTR_PT(334) OR ROM64_INSTR_PT(339)
     OR ROM64_INSTR_PT(340) OR ROM64_INSTR_PT(341)
     OR ROM64_INSTR_PT(342) OR ROM64_INSTR_PT(348)
     OR ROM64_INSTR_PT(350) OR ROM64_INSTR_PT(352)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(359)
     OR ROM64_INSTR_PT(361) OR ROM64_INSTR_PT(364)
     OR ROM64_INSTR_PT(365) OR ROM64_INSTR_PT(366)
     OR ROM64_INSTR_PT(369) OR ROM64_INSTR_PT(371)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(374)
     OR ROM64_INSTR_PT(375) OR ROM64_INSTR_PT(378)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(383) OR ROM64_INSTR_PT(384)
     OR ROM64_INSTR_PT(385) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(389) OR ROM64_INSTR_PT(391)
     OR ROM64_INSTR_PT(394) OR ROM64_INSTR_PT(395)
     OR ROM64_INSTR_PT(396) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(403)
     OR ROM64_INSTR_PT(404) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(406) OR ROM64_INSTR_PT(408)
     OR ROM64_INSTR_PT(409) OR ROM64_INSTR_PT(410)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(419) OR ROM64_INSTR_PT(420)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(424)
     OR ROM64_INSTR_PT(425) OR ROM64_INSTR_PT(426)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(428)
     OR ROM64_INSTR_PT(429) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(437) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(439) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(443)
     OR ROM64_INSTR_PT(445) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(448) OR ROM64_INSTR_PT(451)
     OR ROM64_INSTR_PT(453) OR ROM64_INSTR_PT(454)
     OR ROM64_INSTR_PT(455) OR ROM64_INSTR_PT(456)
     OR ROM64_INSTR_PT(457) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(460) OR ROM64_INSTR_PT(463)
     OR ROM64_INSTR_PT(464) OR ROM64_INSTR_PT(466)
     OR ROM64_INSTR_PT(467) OR ROM64_INSTR_PT(468)
     OR ROM64_INSTR_PT(470) OR ROM64_INSTR_PT(471)
     OR ROM64_INSTR_PT(472) OR ROM64_INSTR_PT(473)
     OR ROM64_INSTR_PT(474) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(478) OR ROM64_INSTR_PT(481)
     OR ROM64_INSTR_PT(482) OR ROM64_INSTR_PT(483)
     OR ROM64_INSTR_PT(484) OR ROM64_INSTR_PT(485)
     OR ROM64_INSTR_PT(488) OR ROM64_INSTR_PT(490)
     OR ROM64_INSTR_PT(491) OR ROM64_INSTR_PT(493)
     OR ROM64_INSTR_PT(495) OR ROM64_INSTR_PT(497)
     OR ROM64_INSTR_PT(498) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(505) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(508) OR ROM64_INSTR_PT(509)
     OR ROM64_INSTR_PT(510) OR ROM64_INSTR_PT(511)
     OR ROM64_INSTR_PT(516) OR ROM64_INSTR_PT(517)
     OR ROM64_INSTR_PT(519) OR ROM64_INSTR_PT(520)
     OR ROM64_INSTR_PT(521) OR ROM64_INSTR_PT(522)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(525)
     OR ROM64_INSTR_PT(532) OR ROM64_INSTR_PT(534)
     OR ROM64_INSTR_PT(538) OR ROM64_INSTR_PT(542)
     OR ROM64_INSTR_PT(546) OR ROM64_INSTR_PT(549)
     OR ROM64_INSTR_PT(551) OR ROM64_INSTR_PT(552)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(555) OR ROM64_INSTR_PT(558)
     OR ROM64_INSTR_PT(559) OR ROM64_INSTR_PT(562)
     OR ROM64_INSTR_PT(563) OR ROM64_INSTR_PT(564)
     OR ROM64_INSTR_PT(566) OR ROM64_INSTR_PT(569)
     OR ROM64_INSTR_PT(570) OR ROM64_INSTR_PT(571)
     OR ROM64_INSTR_PT(572) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(581)
     OR ROM64_INSTR_PT(582) OR ROM64_INSTR_PT(583)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(585)
     OR ROM64_INSTR_PT(586) OR ROM64_INSTR_PT(587)
     OR ROM64_INSTR_PT(588) OR ROM64_INSTR_PT(589)
     OR ROM64_INSTR_PT(590) OR ROM64_INSTR_PT(592)
     OR ROM64_INSTR_PT(595) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(598)
     OR ROM64_INSTR_PT(600) OR ROM64_INSTR_PT(601)
     OR ROM64_INSTR_PT(603) OR ROM64_INSTR_PT(604)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(610) OR ROM64_INSTR_PT(611)
     OR ROM64_INSTR_PT(612) OR ROM64_INSTR_PT(613)
     OR ROM64_INSTR_PT(614) OR ROM64_INSTR_PT(615)
     OR ROM64_INSTR_PT(616) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(620)
     OR ROM64_INSTR_PT(623) OR ROM64_INSTR_PT(626)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(629) OR ROM64_INSTR_PT(632)
     OR ROM64_INSTR_PT(633) OR ROM64_INSTR_PT(635)
     OR ROM64_INSTR_PT(636) OR ROM64_INSTR_PT(639)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(644)
     OR ROM64_INSTR_PT(654) OR ROM64_INSTR_PT(657)
     OR ROM64_INSTR_PT(659) OR ROM64_INSTR_PT(660)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(664)
     OR ROM64_INSTR_PT(666) OR ROM64_INSTR_PT(668)
     OR ROM64_INSTR_PT(675) OR ROM64_INSTR_PT(678)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(682)
     OR ROM64_INSTR_PT(691) OR ROM64_INSTR_PT(695)
     OR ROM64_INSTR_PT(703) OR ROM64_INSTR_PT(706)
     OR ROM64_INSTR_PT(709) OR ROM64_INSTR_PT(713)
     OR ROM64_INSTR_PT(717) OR ROM64_INSTR_PT(721)
     OR ROM64_INSTR_PT(722) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(728)
     OR ROM64_INSTR_PT(731) OR ROM64_INSTR_PT(733)
     OR ROM64_INSTR_PT(735) OR ROM64_INSTR_PT(736)
     OR ROM64_INSTR_PT(738) OR ROM64_INSTR_PT(744)
     OR ROM64_INSTR_PT(759) OR ROM64_INSTR_PT(761)
     OR ROM64_INSTR_PT(766) OR ROM64_INSTR_PT(769)
     OR ROM64_INSTR_PT(776) OR ROM64_INSTR_PT(781)
     OR ROM64_INSTR_PT(794) OR ROM64_INSTR_PT(797)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(809)
     OR ROM64_INSTR_PT(811) OR ROM64_INSTR_PT(813)
     OR ROM64_INSTR_PT(822) OR ROM64_INSTR_PT(824)
     OR ROM64_INSTR_PT(834) OR ROM64_INSTR_PT(846)
     OR ROM64_INSTR_PT(854) OR ROM64_INSTR_PT(855)
     OR ROM64_INSTR_PT(856) OR ROM64_INSTR_PT(858)
     OR ROM64_INSTR_PT(864) OR ROM64_INSTR_PT(869)
     OR ROM64_INSTR_PT(870) OR ROM64_INSTR_PT(883)
    );
MQQ895:TEMPLATE(4) <= 
    (ROM64_INSTR_PT(2) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(10)
     OR ROM64_INSTR_PT(14) OR ROM64_INSTR_PT(15)
     OR ROM64_INSTR_PT(18) OR ROM64_INSTR_PT(20)
     OR ROM64_INSTR_PT(25) OR ROM64_INSTR_PT(28)
     OR ROM64_INSTR_PT(29) OR ROM64_INSTR_PT(33)
     OR ROM64_INSTR_PT(35) OR ROM64_INSTR_PT(36)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(43)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(53)
     OR ROM64_INSTR_PT(56) OR ROM64_INSTR_PT(60)
     OR ROM64_INSTR_PT(65) OR ROM64_INSTR_PT(66)
     OR ROM64_INSTR_PT(69) OR ROM64_INSTR_PT(73)
     OR ROM64_INSTR_PT(74) OR ROM64_INSTR_PT(77)
     OR ROM64_INSTR_PT(78) OR ROM64_INSTR_PT(79)
     OR ROM64_INSTR_PT(80) OR ROM64_INSTR_PT(82)
     OR ROM64_INSTR_PT(84) OR ROM64_INSTR_PT(89)
     OR ROM64_INSTR_PT(92) OR ROM64_INSTR_PT(95)
     OR ROM64_INSTR_PT(96) OR ROM64_INSTR_PT(97)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(101)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(106)
     OR ROM64_INSTR_PT(108) OR ROM64_INSTR_PT(109)
     OR ROM64_INSTR_PT(110) OR ROM64_INSTR_PT(112)
     OR ROM64_INSTR_PT(114) OR ROM64_INSTR_PT(116)
     OR ROM64_INSTR_PT(119) OR ROM64_INSTR_PT(124)
     OR ROM64_INSTR_PT(129) OR ROM64_INSTR_PT(139)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(142)
     OR ROM64_INSTR_PT(143) OR ROM64_INSTR_PT(145)
     OR ROM64_INSTR_PT(146) OR ROM64_INSTR_PT(147)
     OR ROM64_INSTR_PT(150) OR ROM64_INSTR_PT(151)
     OR ROM64_INSTR_PT(153) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(158) OR ROM64_INSTR_PT(160)
     OR ROM64_INSTR_PT(161) OR ROM64_INSTR_PT(166)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(172)
     OR ROM64_INSTR_PT(173) OR ROM64_INSTR_PT(174)
     OR ROM64_INSTR_PT(175) OR ROM64_INSTR_PT(176)
     OR ROM64_INSTR_PT(177) OR ROM64_INSTR_PT(179)
     OR ROM64_INSTR_PT(181) OR ROM64_INSTR_PT(182)
     OR ROM64_INSTR_PT(183) OR ROM64_INSTR_PT(184)
     OR ROM64_INSTR_PT(187) OR ROM64_INSTR_PT(188)
     OR ROM64_INSTR_PT(191) OR ROM64_INSTR_PT(193)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(202)
     OR ROM64_INSTR_PT(203) OR ROM64_INSTR_PT(205)
     OR ROM64_INSTR_PT(206) OR ROM64_INSTR_PT(207)
     OR ROM64_INSTR_PT(208) OR ROM64_INSTR_PT(209)
     OR ROM64_INSTR_PT(211) OR ROM64_INSTR_PT(216)
     OR ROM64_INSTR_PT(219) OR ROM64_INSTR_PT(221)
     OR ROM64_INSTR_PT(225) OR ROM64_INSTR_PT(228)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(231) OR ROM64_INSTR_PT(233)
     OR ROM64_INSTR_PT(237) OR ROM64_INSTR_PT(240)
     OR ROM64_INSTR_PT(242) OR ROM64_INSTR_PT(243)
     OR ROM64_INSTR_PT(247) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(254) OR ROM64_INSTR_PT(257)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(259)
     OR ROM64_INSTR_PT(260) OR ROM64_INSTR_PT(261)
     OR ROM64_INSTR_PT(265) OR ROM64_INSTR_PT(269)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(274)
     OR ROM64_INSTR_PT(277) OR ROM64_INSTR_PT(281)
     OR ROM64_INSTR_PT(284) OR ROM64_INSTR_PT(288)
     OR ROM64_INSTR_PT(290) OR ROM64_INSTR_PT(292)
     OR ROM64_INSTR_PT(294) OR ROM64_INSTR_PT(295)
     OR ROM64_INSTR_PT(304) OR ROM64_INSTR_PT(307)
     OR ROM64_INSTR_PT(309) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(313) OR ROM64_INSTR_PT(319)
     OR ROM64_INSTR_PT(320) OR ROM64_INSTR_PT(324)
     OR ROM64_INSTR_PT(325) OR ROM64_INSTR_PT(327)
     OR ROM64_INSTR_PT(332) OR ROM64_INSTR_PT(334)
     OR ROM64_INSTR_PT(339) OR ROM64_INSTR_PT(340)
     OR ROM64_INSTR_PT(341) OR ROM64_INSTR_PT(342)
     OR ROM64_INSTR_PT(348) OR ROM64_INSTR_PT(350)
     OR ROM64_INSTR_PT(352) OR ROM64_INSTR_PT(353)
     OR ROM64_INSTR_PT(358) OR ROM64_INSTR_PT(359)
     OR ROM64_INSTR_PT(360) OR ROM64_INSTR_PT(361)
     OR ROM64_INSTR_PT(362) OR ROM64_INSTR_PT(365)
     OR ROM64_INSTR_PT(366) OR ROM64_INSTR_PT(368)
     OR ROM64_INSTR_PT(369) OR ROM64_INSTR_PT(371)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(374)
     OR ROM64_INSTR_PT(377) OR ROM64_INSTR_PT(378)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(389) OR ROM64_INSTR_PT(392)
     OR ROM64_INSTR_PT(394) OR ROM64_INSTR_PT(395)
     OR ROM64_INSTR_PT(396) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(402) OR ROM64_INSTR_PT(403)
     OR ROM64_INSTR_PT(405) OR ROM64_INSTR_PT(406)
     OR ROM64_INSTR_PT(408) OR ROM64_INSTR_PT(409)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(419) OR ROM64_INSTR_PT(420)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(425)
     OR ROM64_INSTR_PT(426) OR ROM64_INSTR_PT(428)
     OR ROM64_INSTR_PT(429) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(438) OR ROM64_INSTR_PT(439)
     OR ROM64_INSTR_PT(440) OR ROM64_INSTR_PT(443)
     OR ROM64_INSTR_PT(445) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(448) OR ROM64_INSTR_PT(451)
     OR ROM64_INSTR_PT(453) OR ROM64_INSTR_PT(454)
     OR ROM64_INSTR_PT(455) OR ROM64_INSTR_PT(456)
     OR ROM64_INSTR_PT(458) OR ROM64_INSTR_PT(460)
     OR ROM64_INSTR_PT(463) OR ROM64_INSTR_PT(464)
     OR ROM64_INSTR_PT(466) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(468) OR ROM64_INSTR_PT(470)
     OR ROM64_INSTR_PT(471) OR ROM64_INSTR_PT(472)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(474)
     OR ROM64_INSTR_PT(475) OR ROM64_INSTR_PT(477)
     OR ROM64_INSTR_PT(483) OR ROM64_INSTR_PT(490)
     OR ROM64_INSTR_PT(491) OR ROM64_INSTR_PT(497)
     OR ROM64_INSTR_PT(498) OR ROM64_INSTR_PT(499)
     OR ROM64_INSTR_PT(503) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(508) OR ROM64_INSTR_PT(510)
     OR ROM64_INSTR_PT(516) OR ROM64_INSTR_PT(517)
     OR ROM64_INSTR_PT(519) OR ROM64_INSTR_PT(520)
     OR ROM64_INSTR_PT(527) OR ROM64_INSTR_PT(532)
     OR ROM64_INSTR_PT(538) OR ROM64_INSTR_PT(542)
     OR ROM64_INSTR_PT(546) OR ROM64_INSTR_PT(549)
     OR ROM64_INSTR_PT(551) OR ROM64_INSTR_PT(553)
     OR ROM64_INSTR_PT(554) OR ROM64_INSTR_PT(557)
     OR ROM64_INSTR_PT(559) OR ROM64_INSTR_PT(562)
     OR ROM64_INSTR_PT(564) OR ROM64_INSTR_PT(566)
     OR ROM64_INSTR_PT(570) OR ROM64_INSTR_PT(571)
     OR ROM64_INSTR_PT(572) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(581)
     OR ROM64_INSTR_PT(586) OR ROM64_INSTR_PT(589)
     OR ROM64_INSTR_PT(590) OR ROM64_INSTR_PT(593)
     OR ROM64_INSTR_PT(596) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(598) OR ROM64_INSTR_PT(601)
     OR ROM64_INSTR_PT(602) OR ROM64_INSTR_PT(603)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(606)
     OR ROM64_INSTR_PT(610) OR ROM64_INSTR_PT(611)
     OR ROM64_INSTR_PT(612) OR ROM64_INSTR_PT(613)
     OR ROM64_INSTR_PT(614) OR ROM64_INSTR_PT(615)
     OR ROM64_INSTR_PT(616) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(620) OR ROM64_INSTR_PT(626)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(632) OR ROM64_INSTR_PT(635)
     OR ROM64_INSTR_PT(636) OR ROM64_INSTR_PT(641)
     OR ROM64_INSTR_PT(653) OR ROM64_INSTR_PT(654)
     OR ROM64_INSTR_PT(659) OR ROM64_INSTR_PT(660)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(664)
     OR ROM64_INSTR_PT(668) OR ROM64_INSTR_PT(675)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(682)
     OR ROM64_INSTR_PT(685) OR ROM64_INSTR_PT(691)
     OR ROM64_INSTR_PT(694) OR ROM64_INSTR_PT(695)
     OR ROM64_INSTR_PT(702) OR ROM64_INSTR_PT(703)
     OR ROM64_INSTR_PT(706) OR ROM64_INSTR_PT(709)
     OR ROM64_INSTR_PT(713) OR ROM64_INSTR_PT(716)
     OR ROM64_INSTR_PT(717) OR ROM64_INSTR_PT(721)
     OR ROM64_INSTR_PT(723) OR ROM64_INSTR_PT(724)
     OR ROM64_INSTR_PT(728) OR ROM64_INSTR_PT(733)
     OR ROM64_INSTR_PT(735) OR ROM64_INSTR_PT(736)
     OR ROM64_INSTR_PT(738) OR ROM64_INSTR_PT(741)
     OR ROM64_INSTR_PT(759) OR ROM64_INSTR_PT(766)
     OR ROM64_INSTR_PT(770) OR ROM64_INSTR_PT(781)
     OR ROM64_INSTR_PT(794) OR ROM64_INSTR_PT(797)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(801)
     OR ROM64_INSTR_PT(808) OR ROM64_INSTR_PT(809)
     OR ROM64_INSTR_PT(811) OR ROM64_INSTR_PT(813)
     OR ROM64_INSTR_PT(822) OR ROM64_INSTR_PT(824)
     OR ROM64_INSTR_PT(832) OR ROM64_INSTR_PT(834)
     OR ROM64_INSTR_PT(846) OR ROM64_INSTR_PT(849)
     OR ROM64_INSTR_PT(852) OR ROM64_INSTR_PT(854)
     OR ROM64_INSTR_PT(855) OR ROM64_INSTR_PT(858)
     OR ROM64_INSTR_PT(869) OR ROM64_INSTR_PT(873)
     OR ROM64_INSTR_PT(883));
MQQ896:TEMPLATE(5) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(6)
     OR ROM64_INSTR_PT(7) OR ROM64_INSTR_PT(8)
     OR ROM64_INSTR_PT(11) OR ROM64_INSTR_PT(14)
     OR ROM64_INSTR_PT(15) OR ROM64_INSTR_PT(18)
     OR ROM64_INSTR_PT(21) OR ROM64_INSTR_PT(35)
     OR ROM64_INSTR_PT(38) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(45)
     OR ROM64_INSTR_PT(49) OR ROM64_INSTR_PT(51)
     OR ROM64_INSTR_PT(52) OR ROM64_INSTR_PT(53)
     OR ROM64_INSTR_PT(56) OR ROM64_INSTR_PT(57)
     OR ROM64_INSTR_PT(61) OR ROM64_INSTR_PT(64)
     OR ROM64_INSTR_PT(68) OR ROM64_INSTR_PT(69)
     OR ROM64_INSTR_PT(70) OR ROM64_INSTR_PT(73)
     OR ROM64_INSTR_PT(82) OR ROM64_INSTR_PT(83)
     OR ROM64_INSTR_PT(84) OR ROM64_INSTR_PT(86)
     OR ROM64_INSTR_PT(90) OR ROM64_INSTR_PT(93)
     OR ROM64_INSTR_PT(95) OR ROM64_INSTR_PT(100)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(102)
     OR ROM64_INSTR_PT(105) OR ROM64_INSTR_PT(108)
     OR ROM64_INSTR_PT(109) OR ROM64_INSTR_PT(115)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(124)
     OR ROM64_INSTR_PT(128) OR ROM64_INSTR_PT(132)
     OR ROM64_INSTR_PT(133) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(143)
     OR ROM64_INSTR_PT(144) OR ROM64_INSTR_PT(145)
     OR ROM64_INSTR_PT(153) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(157) OR ROM64_INSTR_PT(158)
     OR ROM64_INSTR_PT(162) OR ROM64_INSTR_PT(164)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(169)
     OR ROM64_INSTR_PT(170) OR ROM64_INSTR_PT(177)
     OR ROM64_INSTR_PT(180) OR ROM64_INSTR_PT(181)
     OR ROM64_INSTR_PT(183) OR ROM64_INSTR_PT(185)
     OR ROM64_INSTR_PT(186) OR ROM64_INSTR_PT(194)
     OR ROM64_INSTR_PT(196) OR ROM64_INSTR_PT(201)
     OR ROM64_INSTR_PT(203) OR ROM64_INSTR_PT(204)
     OR ROM64_INSTR_PT(205) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(211) OR ROM64_INSTR_PT(215)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(219)
     OR ROM64_INSTR_PT(223) OR ROM64_INSTR_PT(226)
     OR ROM64_INSTR_PT(233) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(241) OR ROM64_INSTR_PT(243)
     OR ROM64_INSTR_PT(244) OR ROM64_INSTR_PT(245)
     OR ROM64_INSTR_PT(249) OR ROM64_INSTR_PT(254)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(263) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(265) OR ROM64_INSTR_PT(268)
     OR ROM64_INSTR_PT(269) OR ROM64_INSTR_PT(270)
     OR ROM64_INSTR_PT(272) OR ROM64_INSTR_PT(276)
     OR ROM64_INSTR_PT(278) OR ROM64_INSTR_PT(280)
     OR ROM64_INSTR_PT(282) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(285) OR ROM64_INSTR_PT(287)
     OR ROM64_INSTR_PT(290) OR ROM64_INSTR_PT(293)
     OR ROM64_INSTR_PT(294) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(302) OR ROM64_INSTR_PT(305)
     OR ROM64_INSTR_PT(308) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(312) OR ROM64_INSTR_PT(319)
     OR ROM64_INSTR_PT(325) OR ROM64_INSTR_PT(339)
     OR ROM64_INSTR_PT(348) OR ROM64_INSTR_PT(350)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(355)
     OR ROM64_INSTR_PT(358) OR ROM64_INSTR_PT(364)
     OR ROM64_INSTR_PT(366) OR ROM64_INSTR_PT(367)
     OR ROM64_INSTR_PT(370) OR ROM64_INSTR_PT(372)
     OR ROM64_INSTR_PT(375) OR ROM64_INSTR_PT(378)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(383)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(385)
     OR ROM64_INSTR_PT(391) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(399) OR ROM64_INSTR_PT(403)
     OR ROM64_INSTR_PT(405) OR ROM64_INSTR_PT(409)
     OR ROM64_INSTR_PT(410) OR ROM64_INSTR_PT(413)
     OR ROM64_INSTR_PT(416) OR ROM64_INSTR_PT(417)
     OR ROM64_INSTR_PT(418) OR ROM64_INSTR_PT(419)
     OR ROM64_INSTR_PT(425) OR ROM64_INSTR_PT(426)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(428)
     OR ROM64_INSTR_PT(429) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(432) OR ROM64_INSTR_PT(433)
     OR ROM64_INSTR_PT(435) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(439) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(443)
     OR ROM64_INSTR_PT(445) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(451) OR ROM64_INSTR_PT(453)
     OR ROM64_INSTR_PT(454) OR ROM64_INSTR_PT(455)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(457)
     OR ROM64_INSTR_PT(460) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(478) OR ROM64_INSTR_PT(481)
     OR ROM64_INSTR_PT(482) OR ROM64_INSTR_PT(484)
     OR ROM64_INSTR_PT(485) OR ROM64_INSTR_PT(488)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(493)
     OR ROM64_INSTR_PT(495) OR ROM64_INSTR_PT(496)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(510) OR ROM64_INSTR_PT(512)
     OR ROM64_INSTR_PT(514) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(522) OR ROM64_INSTR_PT(523)
     OR ROM64_INSTR_PT(525) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(531) OR ROM64_INSTR_PT(532)
     OR ROM64_INSTR_PT(534) OR ROM64_INSTR_PT(539)
     OR ROM64_INSTR_PT(542) OR ROM64_INSTR_PT(546)
     OR ROM64_INSTR_PT(552) OR ROM64_INSTR_PT(553)
     OR ROM64_INSTR_PT(554) OR ROM64_INSTR_PT(555)
     OR ROM64_INSTR_PT(557) OR ROM64_INSTR_PT(559)
     OR ROM64_INSTR_PT(563) OR ROM64_INSTR_PT(564)
     OR ROM64_INSTR_PT(566) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(570) OR ROM64_INSTR_PT(571)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(577)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(581)
     OR ROM64_INSTR_PT(582) OR ROM64_INSTR_PT(583)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(585)
     OR ROM64_INSTR_PT(586) OR ROM64_INSTR_PT(587)
     OR ROM64_INSTR_PT(589) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(592) OR ROM64_INSTR_PT(604)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(607)
     OR ROM64_INSTR_PT(608) OR ROM64_INSTR_PT(611)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(616)
     OR ROM64_INSTR_PT(619) OR ROM64_INSTR_PT(625)
     OR ROM64_INSTR_PT(626) OR ROM64_INSTR_PT(627)
     OR ROM64_INSTR_PT(629) OR ROM64_INSTR_PT(633)
     OR ROM64_INSTR_PT(636) OR ROM64_INSTR_PT(639)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(643)
     OR ROM64_INSTR_PT(655) OR ROM64_INSTR_PT(660)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(664)
     OR ROM64_INSTR_PT(666) OR ROM64_INSTR_PT(678)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(695)
     OR ROM64_INSTR_PT(698) OR ROM64_INSTR_PT(702)
     OR ROM64_INSTR_PT(713) OR ROM64_INSTR_PT(716)
     OR ROM64_INSTR_PT(721) OR ROM64_INSTR_PT(722)
     OR ROM64_INSTR_PT(731) OR ROM64_INSTR_PT(736)
     OR ROM64_INSTR_PT(753) OR ROM64_INSTR_PT(761)
     OR ROM64_INSTR_PT(769) OR ROM64_INSTR_PT(770)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(811)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(823)
     OR ROM64_INSTR_PT(824) OR ROM64_INSTR_PT(832)
     OR ROM64_INSTR_PT(834) OR ROM64_INSTR_PT(846)
     OR ROM64_INSTR_PT(854) OR ROM64_INSTR_PT(855)
     OR ROM64_INSTR_PT(856) OR ROM64_INSTR_PT(858)
     OR ROM64_INSTR_PT(864) OR ROM64_INSTR_PT(870)
     OR ROM64_INSTR_PT(873));
MQQ897:TEMPLATE(6) <= 
    ('0');
MQQ898:TEMPLATE(7) <= 
    ('0');
MQQ899:TEMPLATE(8) <= 
    ('0');
MQQ900:TEMPLATE(9) <= 
    (ROM64_INSTR_PT(7) OR ROM64_INSTR_PT(9)
     OR ROM64_INSTR_PT(11) OR ROM64_INSTR_PT(13)
     OR ROM64_INSTR_PT(15) OR ROM64_INSTR_PT(22)
     OR ROM64_INSTR_PT(25) OR ROM64_INSTR_PT(29)
     OR ROM64_INSTR_PT(36) OR ROM64_INSTR_PT(38)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(45)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(55)
     OR ROM64_INSTR_PT(56) OR ROM64_INSTR_PT(58)
     OR ROM64_INSTR_PT(61) OR ROM64_INSTR_PT(70)
     OR ROM64_INSTR_PT(71) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(86) OR ROM64_INSTR_PT(90)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(97)
     OR ROM64_INSTR_PT(100) OR ROM64_INSTR_PT(102)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(105)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(119)
     OR ROM64_INSTR_PT(124) OR ROM64_INSTR_PT(132)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(143) OR ROM64_INSTR_PT(144)
     OR ROM64_INSTR_PT(148) OR ROM64_INSTR_PT(154)
     OR ROM64_INSTR_PT(155) OR ROM64_INSTR_PT(160)
     OR ROM64_INSTR_PT(172) OR ROM64_INSTR_PT(174)
     OR ROM64_INSTR_PT(176) OR ROM64_INSTR_PT(177)
     OR ROM64_INSTR_PT(179) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(181) OR ROM64_INSTR_PT(183)
     OR ROM64_INSTR_PT(186) OR ROM64_INSTR_PT(193)
     OR ROM64_INSTR_PT(201) OR ROM64_INSTR_PT(208)
     OR ROM64_INSTR_PT(213) OR ROM64_INSTR_PT(215)
     OR ROM64_INSTR_PT(216) OR ROM64_INSTR_PT(221)
     OR ROM64_INSTR_PT(222) OR ROM64_INSTR_PT(225)
     OR ROM64_INSTR_PT(226) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(240) OR ROM64_INSTR_PT(242)
     OR ROM64_INSTR_PT(243) OR ROM64_INSTR_PT(245)
     OR ROM64_INSTR_PT(249) OR ROM64_INSTR_PT(259)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(262)
     OR ROM64_INSTR_PT(263) OR ROM64_INSTR_PT(265)
     OR ROM64_INSTR_PT(270) OR ROM64_INSTR_PT(274)
     OR ROM64_INSTR_PT(275) OR ROM64_INSTR_PT(276)
     OR ROM64_INSTR_PT(277) OR ROM64_INSTR_PT(282)
     OR ROM64_INSTR_PT(284) OR ROM64_INSTR_PT(285)
     OR ROM64_INSTR_PT(286) OR ROM64_INSTR_PT(292)
     OR ROM64_INSTR_PT(293) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(299) OR ROM64_INSTR_PT(302)
     OR ROM64_INSTR_PT(305) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(315) OR ROM64_INSTR_PT(319)
     OR ROM64_INSTR_PT(320) OR ROM64_INSTR_PT(322)
     OR ROM64_INSTR_PT(341) OR ROM64_INSTR_PT(349)
     OR ROM64_INSTR_PT(355) OR ROM64_INSTR_PT(359)
     OR ROM64_INSTR_PT(362) OR ROM64_INSTR_PT(365)
     OR ROM64_INSTR_PT(366) OR ROM64_INSTR_PT(369)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(379)
     OR ROM64_INSTR_PT(382) OR ROM64_INSTR_PT(383)
     OR ROM64_INSTR_PT(385) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(389) OR ROM64_INSTR_PT(392)
     OR ROM64_INSTR_PT(394) OR ROM64_INSTR_PT(395)
     OR ROM64_INSTR_PT(396) OR ROM64_INSTR_PT(402)
     OR ROM64_INSTR_PT(403) OR ROM64_INSTR_PT(404)
     OR ROM64_INSTR_PT(405) OR ROM64_INSTR_PT(410)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(415)
     OR ROM64_INSTR_PT(418) OR ROM64_INSTR_PT(425)
     OR ROM64_INSTR_PT(426) OR ROM64_INSTR_PT(429)
     OR ROM64_INSTR_PT(434) OR ROM64_INSTR_PT(435)
     OR ROM64_INSTR_PT(437) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(440) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(451)
     OR ROM64_INSTR_PT(453) OR ROM64_INSTR_PT(456)
     OR ROM64_INSTR_PT(457) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(470) OR ROM64_INSTR_PT(473)
     OR ROM64_INSTR_PT(474) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(478) OR ROM64_INSTR_PT(482)
     OR ROM64_INSTR_PT(485) OR ROM64_INSTR_PT(491)
     OR ROM64_INSTR_PT(493) OR ROM64_INSTR_PT(495)
     OR ROM64_INSTR_PT(498) OR ROM64_INSTR_PT(499)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(505)
     OR ROM64_INSTR_PT(507) OR ROM64_INSTR_PT(509)
     OR ROM64_INSTR_PT(517) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(520) OR ROM64_INSTR_PT(521)
     OR ROM64_INSTR_PT(522) OR ROM64_INSTR_PT(532)
     OR ROM64_INSTR_PT(534) OR ROM64_INSTR_PT(535)
     OR ROM64_INSTR_PT(544) OR ROM64_INSTR_PT(546)
     OR ROM64_INSTR_PT(549) OR ROM64_INSTR_PT(552)
     OR ROM64_INSTR_PT(555) OR ROM64_INSTR_PT(558)
     OR ROM64_INSTR_PT(559) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(569) OR ROM64_INSTR_PT(571)
     OR ROM64_INSTR_PT(572) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(590)
     OR ROM64_INSTR_PT(591) OR ROM64_INSTR_PT(592)
     OR ROM64_INSTR_PT(593) OR ROM64_INSTR_PT(595)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(610) OR ROM64_INSTR_PT(612)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(623)
     OR ROM64_INSTR_PT(628) OR ROM64_INSTR_PT(633)
     OR ROM64_INSTR_PT(639) OR ROM64_INSTR_PT(645)
     OR ROM64_INSTR_PT(646) OR ROM64_INSTR_PT(653)
     OR ROM64_INSTR_PT(659) OR ROM64_INSTR_PT(663)
     OR ROM64_INSTR_PT(666) OR ROM64_INSTR_PT(678)
     OR ROM64_INSTR_PT(691) OR ROM64_INSTR_PT(693)
     OR ROM64_INSTR_PT(703) OR ROM64_INSTR_PT(705)
     OR ROM64_INSTR_PT(741) OR ROM64_INSTR_PT(753)
     OR ROM64_INSTR_PT(797) OR ROM64_INSTR_PT(846)
    );
MQQ901:TEMPLATE(10) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(6)
     OR ROM64_INSTR_PT(7) OR ROM64_INSTR_PT(14)
     OR ROM64_INSTR_PT(15) OR ROM64_INSTR_PT(17)
     OR ROM64_INSTR_PT(20) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(45)
     OR ROM64_INSTR_PT(51) OR ROM64_INSTR_PT(52)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(57)
     OR ROM64_INSTR_PT(73) OR ROM64_INSTR_PT(74)
     OR ROM64_INSTR_PT(75) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(99)
     OR ROM64_INSTR_PT(112) OR ROM64_INSTR_PT(113)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(122) OR ROM64_INSTR_PT(125)
     OR ROM64_INSTR_PT(127) OR ROM64_INSTR_PT(128)
     OR ROM64_INSTR_PT(129) OR ROM64_INSTR_PT(132)
     OR ROM64_INSTR_PT(139) OR ROM64_INSTR_PT(140)
     OR ROM64_INSTR_PT(143) OR ROM64_INSTR_PT(153)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(169)
     OR ROM64_INSTR_PT(171) OR ROM64_INSTR_PT(173)
     OR ROM64_INSTR_PT(174) OR ROM64_INSTR_PT(181)
     OR ROM64_INSTR_PT(183) OR ROM64_INSTR_PT(184)
     OR ROM64_INSTR_PT(185) OR ROM64_INSTR_PT(191)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(199)
     OR ROM64_INSTR_PT(202) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(204) OR ROM64_INSTR_PT(213)
     OR ROM64_INSTR_PT(217) OR ROM64_INSTR_PT(219)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(237) OR ROM64_INSTR_PT(240)
     OR ROM64_INSTR_PT(241) OR ROM64_INSTR_PT(252)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(258)
     OR ROM64_INSTR_PT(260) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(271)
     OR ROM64_INSTR_PT(272) OR ROM64_INSTR_PT(273)
     OR ROM64_INSTR_PT(276) OR ROM64_INSTR_PT(278)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(331)
     OR ROM64_INSTR_PT(339) OR ROM64_INSTR_PT(361)
     OR ROM64_INSTR_PT(364) OR ROM64_INSTR_PT(366)
     OR ROM64_INSTR_PT(367) OR ROM64_INSTR_PT(368)
     OR ROM64_INSTR_PT(374) OR ROM64_INSTR_PT(375)
     OR ROM64_INSTR_PT(377) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(391)
     OR ROM64_INSTR_PT(396) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(403) OR ROM64_INSTR_PT(406)
     OR ROM64_INSTR_PT(408) OR ROM64_INSTR_PT(420)
     OR ROM64_INSTR_PT(424) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(442) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(448) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(472) OR ROM64_INSTR_PT(477)
     OR ROM64_INSTR_PT(480) OR ROM64_INSTR_PT(481)
     OR ROM64_INSTR_PT(483) OR ROM64_INSTR_PT(491)
     OR ROM64_INSTR_PT(503) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(507) OR ROM64_INSTR_PT(508)
     OR ROM64_INSTR_PT(511) OR ROM64_INSTR_PT(512)
     OR ROM64_INSTR_PT(519) OR ROM64_INSTR_PT(525)
     OR ROM64_INSTR_PT(527) OR ROM64_INSTR_PT(531)
     OR ROM64_INSTR_PT(532) OR ROM64_INSTR_PT(538)
     OR ROM64_INSTR_PT(539) OR ROM64_INSTR_PT(545)
     OR ROM64_INSTR_PT(548) OR ROM64_INSTR_PT(553)
     OR ROM64_INSTR_PT(554) OR ROM64_INSTR_PT(557)
     OR ROM64_INSTR_PT(562) OR ROM64_INSTR_PT(563)
     OR ROM64_INSTR_PT(571) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(583) OR ROM64_INSTR_PT(588)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(599)
     OR ROM64_INSTR_PT(600) OR ROM64_INSTR_PT(602)
     OR ROM64_INSTR_PT(603) OR ROM64_INSTR_PT(609)
     OR ROM64_INSTR_PT(614) OR ROM64_INSTR_PT(619)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(629)
     OR ROM64_INSTR_PT(632) OR ROM64_INSTR_PT(636)
     OR ROM64_INSTR_PT(637) OR ROM64_INSTR_PT(641)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(644)
     OR ROM64_INSTR_PT(655) OR ROM64_INSTR_PT(682)
     OR ROM64_INSTR_PT(685) OR ROM64_INSTR_PT(691)
     OR ROM64_INSTR_PT(713) OR ROM64_INSTR_PT(717)
     OR ROM64_INSTR_PT(721) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(728)
     OR ROM64_INSTR_PT(733) OR ROM64_INSTR_PT(735)
     OR ROM64_INSTR_PT(736) OR ROM64_INSTR_PT(738)
     OR ROM64_INSTR_PT(739) OR ROM64_INSTR_PT(761)
     OR ROM64_INSTR_PT(770) OR ROM64_INSTR_PT(824)
     OR ROM64_INSTR_PT(858) OR ROM64_INSTR_PT(873)
    );
MQQ902:TEMPLATE(11) <= 
    ('0');
MQQ903:TEMPLATE(12) <= 
    ('0');
MQQ904:TEMPLATE(13) <= 
    ('0');
MQQ905:TEMPLATE(14) <= 
    (ROM64_INSTR_PT(7) OR ROM64_INSTR_PT(11)
     OR ROM64_INSTR_PT(13) OR ROM64_INSTR_PT(15)
     OR ROM64_INSTR_PT(17) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(25) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(36) OR ROM64_INSTR_PT(38)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(52)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(55)
     OR ROM64_INSTR_PT(56) OR ROM64_INSTR_PT(61)
     OR ROM64_INSTR_PT(64) OR ROM64_INSTR_PT(70)
     OR ROM64_INSTR_PT(73) OR ROM64_INSTR_PT(75)
     OR ROM64_INSTR_PT(77) OR ROM64_INSTR_PT(80)
     OR ROM64_INSTR_PT(84) OR ROM64_INSTR_PT(86)
     OR ROM64_INSTR_PT(89) OR ROM64_INSTR_PT(90)
     OR ROM64_INSTR_PT(92) OR ROM64_INSTR_PT(93)
     OR ROM64_INSTR_PT(96) OR ROM64_INSTR_PT(97)
     OR ROM64_INSTR_PT(99) OR ROM64_INSTR_PT(102)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(106)
     OR ROM64_INSTR_PT(110) OR ROM64_INSTR_PT(113)
     OR ROM64_INSTR_PT(114) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(125)
     OR ROM64_INSTR_PT(127) OR ROM64_INSTR_PT(128)
     OR ROM64_INSTR_PT(132) OR ROM64_INSTR_PT(139)
     OR ROM64_INSTR_PT(144) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(169) OR ROM64_INSTR_PT(171)
     OR ROM64_INSTR_PT(172) OR ROM64_INSTR_PT(174)
     OR ROM64_INSTR_PT(180) OR ROM64_INSTR_PT(181)
     OR ROM64_INSTR_PT(184) OR ROM64_INSTR_PT(186)
     OR ROM64_INSTR_PT(196) OR ROM64_INSTR_PT(199)
     OR ROM64_INSTR_PT(201) OR ROM64_INSTR_PT(202)
     OR ROM64_INSTR_PT(208) OR ROM64_INSTR_PT(213)
     OR ROM64_INSTR_PT(215) OR ROM64_INSTR_PT(216)
     OR ROM64_INSTR_PT(217) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(226) OR ROM64_INSTR_PT(229)
     OR ROM64_INSTR_PT(230) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(240) OR ROM64_INSTR_PT(252)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(270)
     OR ROM64_INSTR_PT(271) OR ROM64_INSTR_PT(272)
     OR ROM64_INSTR_PT(274) OR ROM64_INSTR_PT(275)
     OR ROM64_INSTR_PT(276) OR ROM64_INSTR_PT(277)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(282)
     OR ROM64_INSTR_PT(286) OR ROM64_INSTR_PT(287)
     OR ROM64_INSTR_PT(293) OR ROM64_INSTR_PT(294)
     OR ROM64_INSTR_PT(298) OR ROM64_INSTR_PT(302)
     OR ROM64_INSTR_PT(305) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(315) OR ROM64_INSTR_PT(322)
     OR ROM64_INSTR_PT(331) OR ROM64_INSTR_PT(349)
     OR ROM64_INSTR_PT(364) OR ROM64_INSTR_PT(365)
     OR ROM64_INSTR_PT(366) OR ROM64_INSTR_PT(369)
     OR ROM64_INSTR_PT(371) OR ROM64_INSTR_PT(372)
     OR ROM64_INSTR_PT(375) OR ROM64_INSTR_PT(377)
     OR ROM64_INSTR_PT(383) OR ROM64_INSTR_PT(385)
     OR ROM64_INSTR_PT(388) OR ROM64_INSTR_PT(391)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(396)
     OR ROM64_INSTR_PT(397) OR ROM64_INSTR_PT(403)
     OR ROM64_INSTR_PT(404) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(410) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(420)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(424)
     OR ROM64_INSTR_PT(426) OR ROM64_INSTR_PT(427)
     OR ROM64_INSTR_PT(434) OR ROM64_INSTR_PT(437)
     OR ROM64_INSTR_PT(440) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(457)
     OR ROM64_INSTR_PT(466) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(478) OR ROM64_INSTR_PT(482)
     OR ROM64_INSTR_PT(483) OR ROM64_INSTR_PT(484)
     OR ROM64_INSTR_PT(485) OR ROM64_INSTR_PT(488)
     OR ROM64_INSTR_PT(493) OR ROM64_INSTR_PT(495)
     OR ROM64_INSTR_PT(498) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(505) OR ROM64_INSTR_PT(511)
     OR ROM64_INSTR_PT(517) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(520) OR ROM64_INSTR_PT(521)
     OR ROM64_INSTR_PT(522) OR ROM64_INSTR_PT(523)
     OR ROM64_INSTR_PT(525) OR ROM64_INSTR_PT(532)
     OR ROM64_INSTR_PT(534) OR ROM64_INSTR_PT(535)
     OR ROM64_INSTR_PT(537) OR ROM64_INSTR_PT(539)
     OR ROM64_INSTR_PT(542) OR ROM64_INSTR_PT(544)
     OR ROM64_INSTR_PT(545) OR ROM64_INSTR_PT(548)
     OR ROM64_INSTR_PT(549) OR ROM64_INSTR_PT(552)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(555) OR ROM64_INSTR_PT(558)
     OR ROM64_INSTR_PT(568) OR ROM64_INSTR_PT(569)
     OR ROM64_INSTR_PT(571) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(583) OR ROM64_INSTR_PT(584)
     OR ROM64_INSTR_PT(588) OR ROM64_INSTR_PT(592)
     OR ROM64_INSTR_PT(595) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(600) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(609) OR ROM64_INSTR_PT(612)
     OR ROM64_INSTR_PT(613) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(623)
     OR ROM64_INSTR_PT(628) OR ROM64_INSTR_PT(633)
     OR ROM64_INSTR_PT(636) OR ROM64_INSTR_PT(637)
     OR ROM64_INSTR_PT(639) OR ROM64_INSTR_PT(642)
     OR ROM64_INSTR_PT(644) OR ROM64_INSTR_PT(646)
     OR ROM64_INSTR_PT(649) OR ROM64_INSTR_PT(666)
     OR ROM64_INSTR_PT(678) OR ROM64_INSTR_PT(682)
     OR ROM64_INSTR_PT(691) OR ROM64_INSTR_PT(693)
     OR ROM64_INSTR_PT(703) OR ROM64_INSTR_PT(739)
     OR ROM64_INSTR_PT(744) OR ROM64_INSTR_PT(753)
     OR ROM64_INSTR_PT(761) OR ROM64_INSTR_PT(769)
     OR ROM64_INSTR_PT(776) OR ROM64_INSTR_PT(805)
     OR ROM64_INSTR_PT(823) OR ROM64_INSTR_PT(856)
     OR ROM64_INSTR_PT(864) OR ROM64_INSTR_PT(870)
    );
MQQ906:TEMPLATE(15) <= 
    (ROM64_INSTR_PT(9) OR ROM64_INSTR_PT(15)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(53)
     OR ROM64_INSTR_PT(57) OR ROM64_INSTR_PT(71)
     OR ROM64_INSTR_PT(77) OR ROM64_INSTR_PT(80)
     OR ROM64_INSTR_PT(83) OR ROM64_INSTR_PT(89)
     OR ROM64_INSTR_PT(92) OR ROM64_INSTR_PT(96)
     OR ROM64_INSTR_PT(106) OR ROM64_INSTR_PT(110)
     OR ROM64_INSTR_PT(114) OR ROM64_INSTR_PT(116)
     OR ROM64_INSTR_PT(121) OR ROM64_INSTR_PT(122)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(148)
     OR ROM64_INSTR_PT(158) OR ROM64_INSTR_PT(162)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(170)
     OR ROM64_INSTR_PT(173) OR ROM64_INSTR_PT(174)
     OR ROM64_INSTR_PT(175) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(211) OR ROM64_INSTR_PT(213)
     OR ROM64_INSTR_PT(214) OR ROM64_INSTR_PT(218)
     OR ROM64_INSTR_PT(219) OR ROM64_INSTR_PT(222)
     OR ROM64_INSTR_PT(236) OR ROM64_INSTR_PT(240)
     OR ROM64_INSTR_PT(272) OR ROM64_INSTR_PT(273)
     OR ROM64_INSTR_PT(278) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(294) OR ROM64_INSTR_PT(299)
     OR ROM64_INSTR_PT(311) OR ROM64_INSTR_PT(350)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(358)
     OR ROM64_INSTR_PT(363) OR ROM64_INSTR_PT(370)
     OR ROM64_INSTR_PT(371) OR ROM64_INSTR_PT(396)
     OR ROM64_INSTR_PT(399) OR ROM64_INSTR_PT(408)
     OR ROM64_INSTR_PT(416) OR ROM64_INSTR_PT(417)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(425)
     OR ROM64_INSTR_PT(429) OR ROM64_INSTR_PT(433)
     OR ROM64_INSTR_PT(435) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(442) OR ROM64_INSTR_PT(443)
     OR ROM64_INSTR_PT(451) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(461) OR ROM64_INSTR_PT(466)
     OR ROM64_INSTR_PT(474) OR ROM64_INSTR_PT(480)
     OR ROM64_INSTR_PT(506) OR ROM64_INSTR_PT(508)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(532) OR ROM64_INSTR_PT(537)
     OR ROM64_INSTR_PT(562) OR ROM64_INSTR_PT(564)
     OR ROM64_INSTR_PT(581) OR ROM64_INSTR_PT(582)
     OR ROM64_INSTR_PT(585) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(599) OR ROM64_INSTR_PT(603)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(613)
     OR ROM64_INSTR_PT(614) OR ROM64_INSTR_PT(626)
     OR ROM64_INSTR_PT(659) OR ROM64_INSTR_PT(664)
     OR ROM64_INSTR_PT(691) OR ROM64_INSTR_PT(695)
     OR ROM64_INSTR_PT(716) OR ROM64_INSTR_PT(731)
     OR ROM64_INSTR_PT(832) OR ROM64_INSTR_PT(834)
     OR ROM64_INSTR_PT(846) OR ROM64_INSTR_PT(854)
    );
MQQ907:TEMPLATE(16) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(10)
     OR ROM64_INSTR_PT(17) OR ROM64_INSTR_PT(20)
     OR ROM64_INSTR_PT(21) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(49)
     OR ROM64_INSTR_PT(55) OR ROM64_INSTR_PT(64)
     OR ROM64_INSTR_PT(75) OR ROM64_INSTR_PT(77)
     OR ROM64_INSTR_PT(80) OR ROM64_INSTR_PT(83)
     OR ROM64_INSTR_PT(89) OR ROM64_INSTR_PT(96)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(99)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(106)
     OR ROM64_INSTR_PT(110) OR ROM64_INSTR_PT(113)
     OR ROM64_INSTR_PT(114) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(121)
     OR ROM64_INSTR_PT(127) OR ROM64_INSTR_PT(171)
     OR ROM64_INSTR_PT(175) OR ROM64_INSTR_PT(188)
     OR ROM64_INSTR_PT(191) OR ROM64_INSTR_PT(199)
     OR ROM64_INSTR_PT(208) OR ROM64_INSTR_PT(214)
     OR ROM64_INSTR_PT(217) OR ROM64_INSTR_PT(218)
     OR ROM64_INSTR_PT(223) OR ROM64_INSTR_PT(226)
     OR ROM64_INSTR_PT(252) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(257) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(274)
     OR ROM64_INSTR_PT(275) OR ROM64_INSTR_PT(280)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(286)
     OR ROM64_INSTR_PT(315) OR ROM64_INSTR_PT(322)
     OR ROM64_INSTR_PT(331) OR ROM64_INSTR_PT(349)
     OR ROM64_INSTR_PT(363) OR ROM64_INSTR_PT(369)
     OR ROM64_INSTR_PT(371) OR ROM64_INSTR_PT(375)
     OR ROM64_INSTR_PT(391) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(404)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(422)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(437)
     OR ROM64_INSTR_PT(448) OR ROM64_INSTR_PT(466)
     OR ROM64_INSTR_PT(472) OR ROM64_INSTR_PT(481)
     OR ROM64_INSTR_PT(505) OR ROM64_INSTR_PT(521)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(525)
     OR ROM64_INSTR_PT(538) OR ROM64_INSTR_PT(540)
     OR ROM64_INSTR_PT(558) OR ROM64_INSTR_PT(563)
     OR ROM64_INSTR_PT(569) OR ROM64_INSTR_PT(582)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(595)
     OR ROM64_INSTR_PT(596) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(598) OR ROM64_INSTR_PT(600)
     OR ROM64_INSTR_PT(608) OR ROM64_INSTR_PT(613)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(629)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(644)
     OR ROM64_INSTR_PT(744) OR ROM64_INSTR_PT(769)
     OR ROM64_INSTR_PT(776) OR ROM64_INSTR_PT(870)
    );
MQQ908:TEMPLATE(17) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(17)
     OR ROM64_INSTR_PT(20) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(34) OR ROM64_INSTR_PT(38)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(43)
     OR ROM64_INSTR_PT(49) OR ROM64_INSTR_PT(55)
     OR ROM64_INSTR_PT(61) OR ROM64_INSTR_PT(70)
     OR ROM64_INSTR_PT(77) OR ROM64_INSTR_PT(78)
     OR ROM64_INSTR_PT(80) OR ROM64_INSTR_PT(86)
     OR ROM64_INSTR_PT(89) OR ROM64_INSTR_PT(90)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(99)
     OR ROM64_INSTR_PT(102) OR ROM64_INSTR_PT(104)
     OR ROM64_INSTR_PT(106) OR ROM64_INSTR_PT(111)
     OR ROM64_INSTR_PT(114) OR ROM64_INSTR_PT(118)
     OR ROM64_INSTR_PT(121) OR ROM64_INSTR_PT(127)
     OR ROM64_INSTR_PT(144) OR ROM64_INSTR_PT(168)
     OR ROM64_INSTR_PT(173) OR ROM64_INSTR_PT(175)
     OR ROM64_INSTR_PT(186) OR ROM64_INSTR_PT(188)
     OR ROM64_INSTR_PT(191) OR ROM64_INSTR_PT(199)
     OR ROM64_INSTR_PT(208) OR ROM64_INSTR_PT(215)
     OR ROM64_INSTR_PT(219) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(226) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(252) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(257) OR ROM64_INSTR_PT(270)
     OR ROM64_INSTR_PT(271) OR ROM64_INSTR_PT(274)
     OR ROM64_INSTR_PT(277) OR ROM64_INSTR_PT(280)
     OR ROM64_INSTR_PT(282) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(286) OR ROM64_INSTR_PT(287)
     OR ROM64_INSTR_PT(293) OR ROM64_INSTR_PT(302)
     OR ROM64_INSTR_PT(305) OR ROM64_INSTR_PT(322)
     OR ROM64_INSTR_PT(329) OR ROM64_INSTR_PT(331)
     OR ROM64_INSTR_PT(343) OR ROM64_INSTR_PT(349)
     OR ROM64_INSTR_PT(361) OR ROM64_INSTR_PT(364)
     OR ROM64_INSTR_PT(369) OR ROM64_INSTR_PT(383)
     OR ROM64_INSTR_PT(385) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(406)
     OR ROM64_INSTR_PT(408) OR ROM64_INSTR_PT(410)
     OR ROM64_INSTR_PT(420) OR ROM64_INSTR_PT(422)
     OR ROM64_INSTR_PT(424) OR ROM64_INSTR_PT(427)
     OR ROM64_INSTR_PT(448) OR ROM64_INSTR_PT(466)
     OR ROM64_INSTR_PT(472) OR ROM64_INSTR_PT(478)
     OR ROM64_INSTR_PT(480) OR ROM64_INSTR_PT(481)
     OR ROM64_INSTR_PT(482) OR ROM64_INSTR_PT(483)
     OR ROM64_INSTR_PT(484) OR ROM64_INSTR_PT(485)
     OR ROM64_INSTR_PT(493) OR ROM64_INSTR_PT(495)
     OR ROM64_INSTR_PT(498) OR ROM64_INSTR_PT(508)
     OR ROM64_INSTR_PT(511) OR ROM64_INSTR_PT(522)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(534)
     OR ROM64_INSTR_PT(535) OR ROM64_INSTR_PT(536)
     OR ROM64_INSTR_PT(538) OR ROM64_INSTR_PT(548)
     OR ROM64_INSTR_PT(549) OR ROM64_INSTR_PT(552)
     OR ROM64_INSTR_PT(555) OR ROM64_INSTR_PT(563)
     OR ROM64_INSTR_PT(575) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(583) OR ROM64_INSTR_PT(584)
     OR ROM64_INSTR_PT(588) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(599)
     OR ROM64_INSTR_PT(603) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(612) OR ROM64_INSTR_PT(613)
     OR ROM64_INSTR_PT(614) OR ROM64_INSTR_PT(633)
     OR ROM64_INSTR_PT(637) OR ROM64_INSTR_PT(639)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(644)
     OR ROM64_INSTR_PT(646) OR ROM64_INSTR_PT(666)
     OR ROM64_INSTR_PT(678) OR ROM64_INSTR_PT(682)
     OR ROM64_INSTR_PT(703) OR ROM64_INSTR_PT(870)
    );
MQQ909:TEMPLATE(18) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(20)
     OR ROM64_INSTR_PT(21) OR ROM64_INSTR_PT(39)
     OR ROM64_INSTR_PT(49) OR ROM64_INSTR_PT(77)
     OR ROM64_INSTR_PT(80) OR ROM64_INSTR_PT(89)
     OR ROM64_INSTR_PT(97) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(106) OR ROM64_INSTR_PT(110)
     OR ROM64_INSTR_PT(114) OR ROM64_INSTR_PT(118)
     OR ROM64_INSTR_PT(172) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(273)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(397) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(427)
     OR ROM64_INSTR_PT(466) OR ROM64_INSTR_PT(472)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(538)
     OR ROM64_INSTR_PT(544) OR ROM64_INSTR_PT(563)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(733)
    );
MQQ910:TEMPLATE(19) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(15)
     OR ROM64_INSTR_PT(18) OR ROM64_INSTR_PT(20)
     OR ROM64_INSTR_PT(21) OR ROM64_INSTR_PT(25)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(42)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(49)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(57)
     OR ROM64_INSTR_PT(73) OR ROM64_INSTR_PT(77)
     OR ROM64_INSTR_PT(80) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(97) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(106)
     OR ROM64_INSTR_PT(109) OR ROM64_INSTR_PT(118)
     OR ROM64_INSTR_PT(128) OR ROM64_INSTR_PT(145)
     OR ROM64_INSTR_PT(157) OR ROM64_INSTR_PT(168)
     OR ROM64_INSTR_PT(182) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(205) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(219)
     OR ROM64_INSTR_PT(223) OR ROM64_INSTR_PT(236)
     OR ROM64_INSTR_PT(244) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(254) OR ROM64_INSTR_PT(262)
     OR ROM64_INSTR_PT(269) OR ROM64_INSTR_PT(272)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(280)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(290) OR ROM64_INSTR_PT(308)
     OR ROM64_INSTR_PT(325) OR ROM64_INSTR_PT(348)
     OR ROM64_INSTR_PT(361) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(387) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(397) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(406) OR ROM64_INSTR_PT(409)
     OR ROM64_INSTR_PT(419) OR ROM64_INSTR_PT(422)
     OR ROM64_INSTR_PT(425) OR ROM64_INSTR_PT(427)
     OR ROM64_INSTR_PT(429) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(439) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(451) OR ROM64_INSTR_PT(454)
     OR ROM64_INSTR_PT(455) OR ROM64_INSTR_PT(460)
     OR ROM64_INSTR_PT(466) OR ROM64_INSTR_PT(472)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(510) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(532) OR ROM64_INSTR_PT(538)
     OR ROM64_INSTR_PT(539) OR ROM64_INSTR_PT(542)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(570) OR ROM64_INSTR_PT(577)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(582)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(611) OR ROM64_INSTR_PT(616)
     OR ROM64_INSTR_PT(619) OR ROM64_INSTR_PT(636)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(643)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(733)
     OR ROM64_INSTR_PT(736) OR ROM64_INSTR_PT(770)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(823)
     OR ROM64_INSTR_PT(824));
MQQ911:TEMPLATE(20) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(13)
     OR ROM64_INSTR_PT(18) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(35) OR ROM64_INSTR_PT(36)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(42)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(49)
     OR ROM64_INSTR_PT(56) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(162) OR ROM64_INSTR_PT(196)
     OR ROM64_INSTR_PT(216) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(236) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(262)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(280)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(308) OR ROM64_INSTR_PT(325)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(365)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(425)
     OR ROM64_INSTR_PT(426) OR ROM64_INSTR_PT(427)
     OR ROM64_INSTR_PT(429) OR ROM64_INSTR_PT(435)
     OR ROM64_INSTR_PT(439) OR ROM64_INSTR_PT(451)
     OR ROM64_INSTR_PT(454) OR ROM64_INSTR_PT(455)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(466) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(488) OR ROM64_INSTR_PT(507)
     OR ROM64_INSTR_PT(517) OR ROM64_INSTR_PT(520)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(538)
     OR ROM64_INSTR_PT(542) OR ROM64_INSTR_PT(544)
     OR ROM64_INSTR_PT(564) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(586)
     OR ROM64_INSTR_PT(587) OR ROM64_INSTR_PT(589)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(619) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(681)
     OR ROM64_INSTR_PT(693) OR ROM64_INSTR_PT(721)
     OR ROM64_INSTR_PT(728) OR ROM64_INSTR_PT(735)
     OR ROM64_INSTR_PT(738) OR ROM64_INSTR_PT(770)
     OR ROM64_INSTR_PT(811) OR ROM64_INSTR_PT(823)
    );
MQQ912:TEMPLATE(21) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(6)
     OR ROM64_INSTR_PT(9) OR ROM64_INSTR_PT(10)
     OR ROM64_INSTR_PT(11) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(25)
     OR ROM64_INSTR_PT(36) OR ROM64_INSTR_PT(39)
     OR ROM64_INSTR_PT(43) OR ROM64_INSTR_PT(58)
     OR ROM64_INSTR_PT(70) OR ROM64_INSTR_PT(71)
     OR ROM64_INSTR_PT(76) OR ROM64_INSTR_PT(78)
     OR ROM64_INSTR_PT(83) OR ROM64_INSTR_PT(86)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(96)
     OR ROM64_INSTR_PT(97) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(117) OR ROM64_INSTR_PT(118)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(148)
     OR ROM64_INSTR_PT(154) OR ROM64_INSTR_PT(168)
     OR ROM64_INSTR_PT(172) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(182) OR ROM64_INSTR_PT(184)
     OR ROM64_INSTR_PT(188) OR ROM64_INSTR_PT(194)
     OR ROM64_INSTR_PT(201) OR ROM64_INSTR_PT(202)
     OR ROM64_INSTR_PT(205) OR ROM64_INSTR_PT(214)
     OR ROM64_INSTR_PT(216) OR ROM64_INSTR_PT(219)
     OR ROM64_INSTR_PT(222) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(245) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(257) OR ROM64_INSTR_PT(258)
     OR ROM64_INSTR_PT(260) OR ROM64_INSTR_PT(261)
     OR ROM64_INSTR_PT(264) OR ROM64_INSTR_PT(268)
     OR ROM64_INSTR_PT(271) OR ROM64_INSTR_PT(273)
     OR ROM64_INSTR_PT(275) OR ROM64_INSTR_PT(277)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(298) OR ROM64_INSTR_PT(299)
     OR ROM64_INSTR_PT(312) OR ROM64_INSTR_PT(315)
     OR ROM64_INSTR_PT(348) OR ROM64_INSTR_PT(361)
     OR ROM64_INSTR_PT(363) OR ROM64_INSTR_PT(365)
     OR ROM64_INSTR_PT(371) OR ROM64_INSTR_PT(375)
     OR ROM64_INSTR_PT(387) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(391) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(404)
     OR ROM64_INSTR_PT(406) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(424)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(434) OR ROM64_INSTR_PT(437)
     OR ROM64_INSTR_PT(438) OR ROM64_INSTR_PT(457)
     OR ROM64_INSTR_PT(458) OR ROM64_INSTR_PT(463)
     OR ROM64_INSTR_PT(497) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(505) OR ROM64_INSTR_PT(509)
     OR ROM64_INSTR_PT(510) OR ROM64_INSTR_PT(511)
     OR ROM64_INSTR_PT(520) OR ROM64_INSTR_PT(521)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(525)
     OR ROM64_INSTR_PT(530) OR ROM64_INSTR_PT(531)
     OR ROM64_INSTR_PT(535) OR ROM64_INSTR_PT(538)
     OR ROM64_INSTR_PT(540) OR ROM64_INSTR_PT(544)
     OR ROM64_INSTR_PT(545) OR ROM64_INSTR_PT(549)
     OR ROM64_INSTR_PT(558) OR ROM64_INSTR_PT(569)
     OR ROM64_INSTR_PT(570) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(584)
     OR ROM64_INSTR_PT(588) OR ROM64_INSTR_PT(592)
     OR ROM64_INSTR_PT(595) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(598) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(623)
     OR ROM64_INSTR_PT(628) OR ROM64_INSTR_PT(629)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(728)
     OR ROM64_INSTR_PT(735) OR ROM64_INSTR_PT(738)
     OR ROM64_INSTR_PT(822));
MQQ913:TEMPLATE(22) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(8)
     OR ROM64_INSTR_PT(9) OR ROM64_INSTR_PT(11)
     OR ROM64_INSTR_PT(13) OR ROM64_INSTR_PT(15)
     OR ROM64_INSTR_PT(18) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(25)
     OR ROM64_INSTR_PT(30) OR ROM64_INSTR_PT(36)
     OR ROM64_INSTR_PT(39) OR ROM64_INSTR_PT(43)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(56)
     OR ROM64_INSTR_PT(57) OR ROM64_INSTR_PT(71)
     OR ROM64_INSTR_PT(73) OR ROM64_INSTR_PT(76)
     OR ROM64_INSTR_PT(78) OR ROM64_INSTR_PT(93)
     OR ROM64_INSTR_PT(97) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(113)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(121)
     OR ROM64_INSTR_PT(128) OR ROM64_INSTR_PT(133)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(148)
     OR ROM64_INSTR_PT(155) OR ROM64_INSTR_PT(157)
     OR ROM64_INSTR_PT(162) OR ROM64_INSTR_PT(164)
     OR ROM64_INSTR_PT(171) OR ROM64_INSTR_PT(172)
     OR ROM64_INSTR_PT(175) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(184) OR ROM64_INSTR_PT(188)
     OR ROM64_INSTR_PT(196) OR ROM64_INSTR_PT(201)
     OR ROM64_INSTR_PT(202) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(206) OR ROM64_INSTR_PT(211)
     OR ROM64_INSTR_PT(216) OR ROM64_INSTR_PT(218)
     OR ROM64_INSTR_PT(222) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(244) OR ROM64_INSTR_PT(245)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(257)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(272)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(280)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(298)
     OR ROM64_INSTR_PT(299) OR ROM64_INSTR_PT(312)
     OR ROM64_INSTR_PT(325) OR ROM64_INSTR_PT(353)
     OR ROM64_INSTR_PT(365) OR ROM64_INSTR_PT(372)
     OR ROM64_INSTR_PT(381) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(414) OR ROM64_INSTR_PT(426)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(434)
     OR ROM64_INSTR_PT(438) OR ROM64_INSTR_PT(439)
     OR ROM64_INSTR_PT(440) OR ROM64_INSTR_PT(443)
     OR ROM64_INSTR_PT(454) OR ROM64_INSTR_PT(455)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(457)
     OR ROM64_INSTR_PT(458) OR ROM64_INSTR_PT(460)
     OR ROM64_INSTR_PT(463) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(481) OR ROM64_INSTR_PT(488)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(497)
     OR ROM64_INSTR_PT(503) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(514)
     OR ROM64_INSTR_PT(519) OR ROM64_INSTR_PT(520)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(532)
     OR ROM64_INSTR_PT(538) OR ROM64_INSTR_PT(539)
     OR ROM64_INSTR_PT(540) OR ROM64_INSTR_PT(544)
     OR ROM64_INSTR_PT(545) OR ROM64_INSTR_PT(553)
     OR ROM64_INSTR_PT(554) OR ROM64_INSTR_PT(566)
     OR ROM64_INSTR_PT(568) OR ROM64_INSTR_PT(576)
     OR ROM64_INSTR_PT(581) OR ROM64_INSTR_PT(582)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(586)
     OR ROM64_INSTR_PT(587) OR ROM64_INSTR_PT(589)
     OR ROM64_INSTR_PT(592) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(598)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(607)
     OR ROM64_INSTR_PT(611) OR ROM64_INSTR_PT(613)
     OR ROM64_INSTR_PT(617) OR ROM64_INSTR_PT(625)
     OR ROM64_INSTR_PT(628) OR ROM64_INSTR_PT(636)
     OR ROM64_INSTR_PT(643) OR ROM64_INSTR_PT(655)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(681)
     OR ROM64_INSTR_PT(698) OR ROM64_INSTR_PT(713)
     OR ROM64_INSTR_PT(723) OR ROM64_INSTR_PT(724)
     OR ROM64_INSTR_PT(728) OR ROM64_INSTR_PT(733)
     OR ROM64_INSTR_PT(735) OR ROM64_INSTR_PT(738)
     OR ROM64_INSTR_PT(822) OR ROM64_INSTR_PT(824)
     OR ROM64_INSTR_PT(846) OR ROM64_INSTR_PT(854)
    );
MQQ914:TEMPLATE(23) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(6)
     OR ROM64_INSTR_PT(13) OR ROM64_INSTR_PT(25)
     OR ROM64_INSTR_PT(36) OR ROM64_INSTR_PT(39)
     OR ROM64_INSTR_PT(56) OR ROM64_INSTR_PT(57)
     OR ROM64_INSTR_PT(73) OR ROM64_INSTR_PT(89)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(100) OR ROM64_INSTR_PT(101)
     OR ROM64_INSTR_PT(110) OR ROM64_INSTR_PT(114)
     OR ROM64_INSTR_PT(124) OR ROM64_INSTR_PT(128)
     OR ROM64_INSTR_PT(137) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(157) OR ROM64_INSTR_PT(162)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(184) OR ROM64_INSTR_PT(194)
     OR ROM64_INSTR_PT(201) OR ROM64_INSTR_PT(202)
     OR ROM64_INSTR_PT(203) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(216) OR ROM64_INSTR_PT(218)
     OR ROM64_INSTR_PT(219) OR ROM64_INSTR_PT(229)
     OR ROM64_INSTR_PT(230) OR ROM64_INSTR_PT(244)
     OR ROM64_INSTR_PT(245) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(263)
     OR ROM64_INSTR_PT(277) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(285) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(312) OR ROM64_INSTR_PT(319)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(361)
     OR ROM64_INSTR_PT(365) OR ROM64_INSTR_PT(372)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(388) OR ROM64_INSTR_PT(395)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(406) OR ROM64_INSTR_PT(413)
     OR ROM64_INSTR_PT(426) OR ROM64_INSTR_PT(434)
     OR ROM64_INSTR_PT(438) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(457)
     OR ROM64_INSTR_PT(458) OR ROM64_INSTR_PT(460)
     OR ROM64_INSTR_PT(467) OR ROM64_INSTR_PT(473)
     OR ROM64_INSTR_PT(475) OR ROM64_INSTR_PT(488)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(517) OR ROM64_INSTR_PT(520)
     OR ROM64_INSTR_PT(531) OR ROM64_INSTR_PT(535)
     OR ROM64_INSTR_PT(538) OR ROM64_INSTR_PT(539)
     OR ROM64_INSTR_PT(545) OR ROM64_INSTR_PT(546)
     OR ROM64_INSTR_PT(549) OR ROM64_INSTR_PT(553)
     OR ROM64_INSTR_PT(554) OR ROM64_INSTR_PT(559)
     OR ROM64_INSTR_PT(563) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(575) OR ROM64_INSTR_PT(582)
     OR ROM64_INSTR_PT(592) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(611)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(623) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(636) OR ROM64_INSTR_PT(643)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(693)
     OR ROM64_INSTR_PT(717) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(728)
     OR ROM64_INSTR_PT(733) OR ROM64_INSTR_PT(735)
     OR ROM64_INSTR_PT(738) OR ROM64_INSTR_PT(822)
     OR ROM64_INSTR_PT(824) OR ROM64_INSTR_PT(846)
    );
MQQ915:TEMPLATE(24) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(11)
     OR ROM64_INSTR_PT(14) OR ROM64_INSTR_PT(30)
     OR ROM64_INSTR_PT(36) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(51)
     OR ROM64_INSTR_PT(77) OR ROM64_INSTR_PT(80)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(100) OR ROM64_INSTR_PT(105)
     OR ROM64_INSTR_PT(106) OR ROM64_INSTR_PT(115)
     OR ROM64_INSTR_PT(124) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(143)
     OR ROM64_INSTR_PT(153) OR ROM64_INSTR_PT(158)
     OR ROM64_INSTR_PT(170) OR ROM64_INSTR_PT(172)
     OR ROM64_INSTR_PT(184) OR ROM64_INSTR_PT(185)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(202)
     OR ROM64_INSTR_PT(204) OR ROM64_INSTR_PT(216)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(229)
     OR ROM64_INSTR_PT(230) OR ROM64_INSTR_PT(241)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(258)
     OR ROM64_INSTR_PT(260) OR ROM64_INSTR_PT(261)
     OR ROM64_INSTR_PT(262) OR ROM64_INSTR_PT(263)
     OR ROM64_INSTR_PT(277) OR ROM64_INSTR_PT(278)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(285)
     OR ROM64_INSTR_PT(294) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(308) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(319) OR ROM64_INSTR_PT(348)
     OR ROM64_INSTR_PT(365) OR ROM64_INSTR_PT(366)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(387)
     OR ROM64_INSTR_PT(394) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(428) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(432) OR ROM64_INSTR_PT(433)
     OR ROM64_INSTR_PT(434) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(453) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(496) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(512)
     OR ROM64_INSTR_PT(520) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(531) OR ROM64_INSTR_PT(535)
     OR ROM64_INSTR_PT(544) OR ROM64_INSTR_PT(545)
     OR ROM64_INSTR_PT(546) OR ROM64_INSTR_PT(549)
     OR ROM64_INSTR_PT(557) OR ROM64_INSTR_PT(559)
     OR ROM64_INSTR_PT(564) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(580)
     OR ROM64_INSTR_PT(582) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(606)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(617)
     OR ROM64_INSTR_PT(619) OR ROM64_INSTR_PT(623)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(645) OR ROM64_INSTR_PT(663)
     OR ROM64_INSTR_PT(693) OR ROM64_INSTR_PT(705)
     OR ROM64_INSTR_PT(736) OR ROM64_INSTR_PT(753)
     OR ROM64_INSTR_PT(770) OR ROM64_INSTR_PT(822)
     OR ROM64_INSTR_PT(846));
MQQ916:TEMPLATE(25) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(6)
     OR ROM64_INSTR_PT(13) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(25) OR ROM64_INSTR_PT(36)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(56)
     OR ROM64_INSTR_PT(57) OR ROM64_INSTR_PT(73)
     OR ROM64_INSTR_PT(97) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(118)
     OR ROM64_INSTR_PT(125) OR ROM64_INSTR_PT(128)
     OR ROM64_INSTR_PT(134) OR ROM64_INSTR_PT(143)
     OR ROM64_INSTR_PT(155) OR ROM64_INSTR_PT(157)
     OR ROM64_INSTR_PT(158) OR ROM64_INSTR_PT(162)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(170)
     OR ROM64_INSTR_PT(172) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(182) OR ROM64_INSTR_PT(184)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(196)
     OR ROM64_INSTR_PT(202) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(206) OR ROM64_INSTR_PT(216)
     OR ROM64_INSTR_PT(219) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(244) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(260) OR ROM64_INSTR_PT(261)
     OR ROM64_INSTR_PT(277) OR ROM64_INSTR_PT(278)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(294) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(339) OR ROM64_INSTR_PT(348)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(361)
     OR ROM64_INSTR_PT(365) OR ROM64_INSTR_PT(366)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(387) OR ROM64_INSTR_PT(395)
     OR ROM64_INSTR_PT(397) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(405) OR ROM64_INSTR_PT(406)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(426)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(433) OR ROM64_INSTR_PT(434)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(460) OR ROM64_INSTR_PT(466)
     OR ROM64_INSTR_PT(467) OR ROM64_INSTR_PT(473)
     OR ROM64_INSTR_PT(475) OR ROM64_INSTR_PT(488)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(506) OR ROM64_INSTR_PT(507)
     OR ROM64_INSTR_PT(517) OR ROM64_INSTR_PT(520)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(531) OR ROM64_INSTR_PT(535)
     OR ROM64_INSTR_PT(539) OR ROM64_INSTR_PT(542)
     OR ROM64_INSTR_PT(545) OR ROM64_INSTR_PT(549)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(557) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(575) OR ROM64_INSTR_PT(576)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(584)
     OR ROM64_INSTR_PT(585) OR ROM64_INSTR_PT(592)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(611)
     OR ROM64_INSTR_PT(617) OR ROM64_INSTR_PT(626)
     OR ROM64_INSTR_PT(632) OR ROM64_INSTR_PT(636)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(643)
     OR ROM64_INSTR_PT(649) OR ROM64_INSTR_PT(655)
     OR ROM64_INSTR_PT(664) OR ROM64_INSTR_PT(693)
     OR ROM64_INSTR_PT(702) OR ROM64_INSTR_PT(713)
     OR ROM64_INSTR_PT(736) OR ROM64_INSTR_PT(739)
     OR ROM64_INSTR_PT(753) OR ROM64_INSTR_PT(798)
     OR ROM64_INSTR_PT(822) OR ROM64_INSTR_PT(823)
     OR ROM64_INSTR_PT(824) OR ROM64_INSTR_PT(832)
    );
MQQ917:TEMPLATE(26) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(7)
     OR ROM64_INSTR_PT(9) OR ROM64_INSTR_PT(11)
     OR ROM64_INSTR_PT(14) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(25)
     OR ROM64_INSTR_PT(30) OR ROM64_INSTR_PT(35)
     OR ROM64_INSTR_PT(36) OR ROM64_INSTR_PT(38)
     OR ROM64_INSTR_PT(41) OR ROM64_INSTR_PT(43)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(50)
     OR ROM64_INSTR_PT(51) OR ROM64_INSTR_PT(52)
     OR ROM64_INSTR_PT(56) OR ROM64_INSTR_PT(57)
     OR ROM64_INSTR_PT(58) OR ROM64_INSTR_PT(61)
     OR ROM64_INSTR_PT(68) OR ROM64_INSTR_PT(69)
     OR ROM64_INSTR_PT(70) OR ROM64_INSTR_PT(71)
     OR ROM64_INSTR_PT(73) OR ROM64_INSTR_PT(76)
     OR ROM64_INSTR_PT(78) OR ROM64_INSTR_PT(82)
     OR ROM64_INSTR_PT(83) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(86) OR ROM64_INSTR_PT(90)
     OR ROM64_INSTR_PT(92) OR ROM64_INSTR_PT(93)
     OR ROM64_INSTR_PT(95) OR ROM64_INSTR_PT(97)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(100)
     OR ROM64_INSTR_PT(101) OR ROM64_INSTR_PT(102)
     OR ROM64_INSTR_PT(105) OR ROM64_INSTR_PT(108)
     OR ROM64_INSTR_PT(109) OR ROM64_INSTR_PT(115)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(124)
     OR ROM64_INSTR_PT(128) OR ROM64_INSTR_PT(132)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(143)
     OR ROM64_INSTR_PT(144) OR ROM64_INSTR_PT(145)
     OR ROM64_INSTR_PT(148) OR ROM64_INSTR_PT(153)
     OR ROM64_INSTR_PT(154) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(157) OR ROM64_INSTR_PT(158)
     OR ROM64_INSTR_PT(162) OR ROM64_INSTR_PT(169)
     OR ROM64_INSTR_PT(172) OR ROM64_INSTR_PT(174)
     OR ROM64_INSTR_PT(177) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(181) OR ROM64_INSTR_PT(183)
     OR ROM64_INSTR_PT(185) OR ROM64_INSTR_PT(186)
     OR ROM64_INSTR_PT(188) OR ROM64_INSTR_PT(194)
     OR ROM64_INSTR_PT(196) OR ROM64_INSTR_PT(201)
     OR ROM64_INSTR_PT(203) OR ROM64_INSTR_PT(204)
     OR ROM64_INSTR_PT(205) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(215) OR ROM64_INSTR_PT(216)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(222)
     OR ROM64_INSTR_PT(223) OR ROM64_INSTR_PT(226)
     OR ROM64_INSTR_PT(233) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(241) OR ROM64_INSTR_PT(243)
     OR ROM64_INSTR_PT(244) OR ROM64_INSTR_PT(245)
     OR ROM64_INSTR_PT(249) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(254) OR ROM64_INSTR_PT(257)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(261) OR ROM64_INSTR_PT(263)
     OR ROM64_INSTR_PT(264) OR ROM64_INSTR_PT(265)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(269)
     OR ROM64_INSTR_PT(270) OR ROM64_INSTR_PT(271)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(275)
     OR ROM64_INSTR_PT(276) OR ROM64_INSTR_PT(277)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(282)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(285) OR ROM64_INSTR_PT(287)
     OR ROM64_INSTR_PT(290) OR ROM64_INSTR_PT(293)
     OR ROM64_INSTR_PT(294) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(298) OR ROM64_INSTR_PT(299)
     OR ROM64_INSTR_PT(302) OR ROM64_INSTR_PT(305)
     OR ROM64_INSTR_PT(308) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(312) OR ROM64_INSTR_PT(315)
     OR ROM64_INSTR_PT(319) OR ROM64_INSTR_PT(339)
     OR ROM64_INSTR_PT(348) OR ROM64_INSTR_PT(350)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(355)
     OR ROM64_INSTR_PT(358) OR ROM64_INSTR_PT(364)
     OR ROM64_INSTR_PT(365) OR ROM64_INSTR_PT(367)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(374)
     OR ROM64_INSTR_PT(375) OR ROM64_INSTR_PT(378)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(383) OR ROM64_INSTR_PT(384)
     OR ROM64_INSTR_PT(385) OR ROM64_INSTR_PT(388)
     OR ROM64_INSTR_PT(391) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(397)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(403)
     OR ROM64_INSTR_PT(404) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(409) OR ROM64_INSTR_PT(410)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(419) OR ROM64_INSTR_PT(424)
     OR ROM64_INSTR_PT(425) OR ROM64_INSTR_PT(426)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(428)
     OR ROM64_INSTR_PT(429) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(432) OR ROM64_INSTR_PT(435)
     OR ROM64_INSTR_PT(437) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(451)
     OR ROM64_INSTR_PT(453) OR ROM64_INSTR_PT(456)
     OR ROM64_INSTR_PT(457) OR ROM64_INSTR_PT(458)
     OR ROM64_INSTR_PT(460) OR ROM64_INSTR_PT(461)
     OR ROM64_INSTR_PT(463) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(478) OR ROM64_INSTR_PT(481)
     OR ROM64_INSTR_PT(482) OR ROM64_INSTR_PT(484)
     OR ROM64_INSTR_PT(485) OR ROM64_INSTR_PT(488)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(493)
     OR ROM64_INSTR_PT(495) OR ROM64_INSTR_PT(496)
     OR ROM64_INSTR_PT(497) OR ROM64_INSTR_PT(504)
     OR ROM64_INSTR_PT(505) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(510)
     OR ROM64_INSTR_PT(511) OR ROM64_INSTR_PT(512)
     OR ROM64_INSTR_PT(517) OR ROM64_INSTR_PT(520)
     OR ROM64_INSTR_PT(521) OR ROM64_INSTR_PT(522)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(525)
     OR ROM64_INSTR_PT(530) OR ROM64_INSTR_PT(531)
     OR ROM64_INSTR_PT(534) OR ROM64_INSTR_PT(535)
     OR ROM64_INSTR_PT(539) OR ROM64_INSTR_PT(540)
     OR ROM64_INSTR_PT(544) OR ROM64_INSTR_PT(546)
     OR ROM64_INSTR_PT(549) OR ROM64_INSTR_PT(552)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(555) OR ROM64_INSTR_PT(557)
     OR ROM64_INSTR_PT(558) OR ROM64_INSTR_PT(559)
     OR ROM64_INSTR_PT(563) OR ROM64_INSTR_PT(564)
     OR ROM64_INSTR_PT(568) OR ROM64_INSTR_PT(569)
     OR ROM64_INSTR_PT(570) OR ROM64_INSTR_PT(571)
     OR ROM64_INSTR_PT(575) OR ROM64_INSTR_PT(576)
     OR ROM64_INSTR_PT(577) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(582)
     OR ROM64_INSTR_PT(583) OR ROM64_INSTR_PT(584)
     OR ROM64_INSTR_PT(588) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(592) OR ROM64_INSTR_PT(595)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(598)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(609) OR ROM64_INSTR_PT(611)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(616)
     OR ROM64_INSTR_PT(617) OR ROM64_INSTR_PT(618)
     OR ROM64_INSTR_PT(619) OR ROM64_INSTR_PT(623)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(629) OR ROM64_INSTR_PT(632)
     OR ROM64_INSTR_PT(633) OR ROM64_INSTR_PT(636)
     OR ROM64_INSTR_PT(639) OR ROM64_INSTR_PT(642)
     OR ROM64_INSTR_PT(643) OR ROM64_INSTR_PT(655)
     OR ROM64_INSTR_PT(660) OR ROM64_INSTR_PT(663)
     OR ROM64_INSTR_PT(664) OR ROM64_INSTR_PT(666)
     OR ROM64_INSTR_PT(678) OR ROM64_INSTR_PT(695)
     OR ROM64_INSTR_PT(702) OR ROM64_INSTR_PT(713)
     OR ROM64_INSTR_PT(716) OR ROM64_INSTR_PT(717)
     OR ROM64_INSTR_PT(721) OR ROM64_INSTR_PT(722)
     OR ROM64_INSTR_PT(723) OR ROM64_INSTR_PT(724)
     OR ROM64_INSTR_PT(733) OR ROM64_INSTR_PT(736)
     OR ROM64_INSTR_PT(761) OR ROM64_INSTR_PT(770)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(811)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(822)
     OR ROM64_INSTR_PT(824) OR ROM64_INSTR_PT(832)
     OR ROM64_INSTR_PT(834) OR ROM64_INSTR_PT(846)
     OR ROM64_INSTR_PT(855) OR ROM64_INSTR_PT(856)
     OR ROM64_INSTR_PT(858) OR ROM64_INSTR_PT(864)
     OR ROM64_INSTR_PT(870) OR ROM64_INSTR_PT(873)
    );
MQQ918:TEMPLATE(27) <= 
    (ROM64_INSTR_PT(5) OR ROM64_INSTR_PT(6)
     OR ROM64_INSTR_PT(7) OR ROM64_INSTR_PT(8)
     OR ROM64_INSTR_PT(9) OR ROM64_INSTR_PT(11)
     OR ROM64_INSTR_PT(15) OR ROM64_INSTR_PT(18)
     OR ROM64_INSTR_PT(21) OR ROM64_INSTR_PT(22)
     OR ROM64_INSTR_PT(35) OR ROM64_INSTR_PT(38)
     OR ROM64_INSTR_PT(42) OR ROM64_INSTR_PT(45)
     OR ROM64_INSTR_PT(49) OR ROM64_INSTR_PT(52)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(56)
     OR ROM64_INSTR_PT(57) OR ROM64_INSTR_PT(61)
     OR ROM64_INSTR_PT(68) OR ROM64_INSTR_PT(69)
     OR ROM64_INSTR_PT(71) OR ROM64_INSTR_PT(73)
     OR ROM64_INSTR_PT(82) OR ROM64_INSTR_PT(83)
     OR ROM64_INSTR_PT(84) OR ROM64_INSTR_PT(90)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(95)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(101)
     OR ROM64_INSTR_PT(102) OR ROM64_INSTR_PT(108)
     OR ROM64_INSTR_PT(109) OR ROM64_INSTR_PT(113)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(118) OR ROM64_INSTR_PT(128)
     OR ROM64_INSTR_PT(132) OR ROM64_INSTR_PT(133)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(143)
     OR ROM64_INSTR_PT(144) OR ROM64_INSTR_PT(145)
     OR ROM64_INSTR_PT(148) OR ROM64_INSTR_PT(155)
     OR ROM64_INSTR_PT(157) OR ROM64_INSTR_PT(158)
     OR ROM64_INSTR_PT(162) OR ROM64_INSTR_PT(164)
     OR ROM64_INSTR_PT(168) OR ROM64_INSTR_PT(169)
     OR ROM64_INSTR_PT(170) OR ROM64_INSTR_PT(171)
     OR ROM64_INSTR_PT(177) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(181) OR ROM64_INSTR_PT(182)
     OR ROM64_INSTR_PT(183) OR ROM64_INSTR_PT(186)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(196)
     OR ROM64_INSTR_PT(201) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(205) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(211) OR ROM64_INSTR_PT(215)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(219)
     OR ROM64_INSTR_PT(222) OR ROM64_INSTR_PT(223)
     OR ROM64_INSTR_PT(226) OR ROM64_INSTR_PT(233)
     OR ROM64_INSTR_PT(238) OR ROM64_INSTR_PT(240)
     OR ROM64_INSTR_PT(243) OR ROM64_INSTR_PT(244)
     OR ROM64_INSTR_PT(245) OR ROM64_INSTR_PT(249)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(254)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(264) OR ROM64_INSTR_PT(265)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(269)
     OR ROM64_INSTR_PT(270) OR ROM64_INSTR_PT(272)
     OR ROM64_INSTR_PT(276) OR ROM64_INSTR_PT(278)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(282)
     OR ROM64_INSTR_PT(283) OR ROM64_INSTR_PT(284)
     OR ROM64_INSTR_PT(287) OR ROM64_INSTR_PT(290)
     OR ROM64_INSTR_PT(293) OR ROM64_INSTR_PT(294)
     OR ROM64_INSTR_PT(298) OR ROM64_INSTR_PT(299)
     OR ROM64_INSTR_PT(302) OR ROM64_INSTR_PT(311)
     OR ROM64_INSTR_PT(312) OR ROM64_INSTR_PT(325)
     OR ROM64_INSTR_PT(339) OR ROM64_INSTR_PT(348)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(361)
     OR ROM64_INSTR_PT(364) OR ROM64_INSTR_PT(366)
     OR ROM64_INSTR_PT(367) OR ROM64_INSTR_PT(372)
     OR ROM64_INSTR_PT(374) OR ROM64_INSTR_PT(375)
     OR ROM64_INSTR_PT(378) OR ROM64_INSTR_PT(381)
     OR ROM64_INSTR_PT(383) OR ROM64_INSTR_PT(384)
     OR ROM64_INSTR_PT(385) OR ROM64_INSTR_PT(391)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(396)
     OR ROM64_INSTR_PT(397) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(403) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(406) OR ROM64_INSTR_PT(409)
     OR ROM64_INSTR_PT(410) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(419) OR ROM64_INSTR_PT(425)
     OR ROM64_INSTR_PT(426) OR ROM64_INSTR_PT(427)
     OR ROM64_INSTR_PT(428) OR ROM64_INSTR_PT(429)
     OR ROM64_INSTR_PT(430) OR ROM64_INSTR_PT(433)
     OR ROM64_INSTR_PT(435) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(439) OR ROM64_INSTR_PT(440)
     OR ROM64_INSTR_PT(443) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(451) OR ROM64_INSTR_PT(454)
     OR ROM64_INSTR_PT(455) OR ROM64_INSTR_PT(456)
     OR ROM64_INSTR_PT(457) OR ROM64_INSTR_PT(460)
     OR ROM64_INSTR_PT(467) OR ROM64_INSTR_PT(473)
     OR ROM64_INSTR_PT(475) OR ROM64_INSTR_PT(478)
     OR ROM64_INSTR_PT(481) OR ROM64_INSTR_PT(482)
     OR ROM64_INSTR_PT(484) OR ROM64_INSTR_PT(485)
     OR ROM64_INSTR_PT(488) OR ROM64_INSTR_PT(490)
     OR ROM64_INSTR_PT(495) OR ROM64_INSTR_PT(506)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(510)
     OR ROM64_INSTR_PT(514) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(522) OR ROM64_INSTR_PT(523)
     OR ROM64_INSTR_PT(525) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(531) OR ROM64_INSTR_PT(532)
     OR ROM64_INSTR_PT(534) OR ROM64_INSTR_PT(539)
     OR ROM64_INSTR_PT(542) OR ROM64_INSTR_PT(552)
     OR ROM64_INSTR_PT(553) OR ROM64_INSTR_PT(554)
     OR ROM64_INSTR_PT(555) OR ROM64_INSTR_PT(557)
     OR ROM64_INSTR_PT(563) OR ROM64_INSTR_PT(564)
     OR ROM64_INSTR_PT(566) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(570) OR ROM64_INSTR_PT(571)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(577)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(581)
     OR ROM64_INSTR_PT(582) OR ROM64_INSTR_PT(583)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(585)
     OR ROM64_INSTR_PT(586) OR ROM64_INSTR_PT(587)
     OR ROM64_INSTR_PT(589) OR ROM64_INSTR_PT(592)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(604)
     OR ROM64_INSTR_PT(607) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(611) OR ROM64_INSTR_PT(616)
     OR ROM64_INSTR_PT(619) OR ROM64_INSTR_PT(625)
     OR ROM64_INSTR_PT(626) OR ROM64_INSTR_PT(629)
     OR ROM64_INSTR_PT(632) OR ROM64_INSTR_PT(633)
     OR ROM64_INSTR_PT(636) OR ROM64_INSTR_PT(639)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(643)
     OR ROM64_INSTR_PT(655) OR ROM64_INSTR_PT(660)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(664)
     OR ROM64_INSTR_PT(666) OR ROM64_INSTR_PT(678)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(698)
     OR ROM64_INSTR_PT(702) OR ROM64_INSTR_PT(713)
     OR ROM64_INSTR_PT(722) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(733)
     OR ROM64_INSTR_PT(736) OR ROM64_INSTR_PT(753)
     OR ROM64_INSTR_PT(761) OR ROM64_INSTR_PT(770)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(811)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(823)
     OR ROM64_INSTR_PT(824) OR ROM64_INSTR_PT(832)
     OR ROM64_INSTR_PT(834) OR ROM64_INSTR_PT(854)
     OR ROM64_INSTR_PT(855) OR ROM64_INSTR_PT(856)
     OR ROM64_INSTR_PT(864) OR ROM64_INSTR_PT(870)
    );
MQQ919:TEMPLATE(28) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(9)
     OR ROM64_INSTR_PT(14) OR ROM64_INSTR_PT(17)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(38) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(51)
     OR ROM64_INSTR_PT(52) OR ROM64_INSTR_PT(56)
     OR ROM64_INSTR_PT(57) OR ROM64_INSTR_PT(61)
     OR ROM64_INSTR_PT(64) OR ROM64_INSTR_PT(68)
     OR ROM64_INSTR_PT(69) OR ROM64_INSTR_PT(70)
     OR ROM64_INSTR_PT(71) OR ROM64_INSTR_PT(73)
     OR ROM64_INSTR_PT(75) OR ROM64_INSTR_PT(82)
     OR ROM64_INSTR_PT(83) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(86) OR ROM64_INSTR_PT(90)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(95)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(99)
     OR ROM64_INSTR_PT(100) OR ROM64_INSTR_PT(101)
     OR ROM64_INSTR_PT(102) OR ROM64_INSTR_PT(105)
     OR ROM64_INSTR_PT(108) OR ROM64_INSTR_PT(113)
     OR ROM64_INSTR_PT(115) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(124) OR ROM64_INSTR_PT(125)
     OR ROM64_INSTR_PT(127) OR ROM64_INSTR_PT(128)
     OR ROM64_INSTR_PT(134) OR ROM64_INSTR_PT(136)
     OR ROM64_INSTR_PT(137) OR ROM64_INSTR_PT(140)
     OR ROM64_INSTR_PT(143) OR ROM64_INSTR_PT(144)
     OR ROM64_INSTR_PT(148) OR ROM64_INSTR_PT(153)
     OR ROM64_INSTR_PT(155) OR ROM64_INSTR_PT(157)
     OR ROM64_INSTR_PT(158) OR ROM64_INSTR_PT(162)
     OR ROM64_INSTR_PT(169) OR ROM64_INSTR_PT(171)
     OR ROM64_INSTR_PT(180) OR ROM64_INSTR_PT(185)
     OR ROM64_INSTR_PT(186) OR ROM64_INSTR_PT(194)
     OR ROM64_INSTR_PT(196) OR ROM64_INSTR_PT(199)
     OR ROM64_INSTR_PT(201) OR ROM64_INSTR_PT(203)
     OR ROM64_INSTR_PT(204) OR ROM64_INSTR_PT(206)
     OR ROM64_INSTR_PT(215) OR ROM64_INSTR_PT(217)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(222)
     OR ROM64_INSTR_PT(226) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(241) OR ROM64_INSTR_PT(243)
     OR ROM64_INSTR_PT(244) OR ROM64_INSTR_PT(249)
     OR ROM64_INSTR_PT(252) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(263) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(265) OR ROM64_INSTR_PT(268)
     OR ROM64_INSTR_PT(269) OR ROM64_INSTR_PT(270)
     OR ROM64_INSTR_PT(271) OR ROM64_INSTR_PT(275)
     OR ROM64_INSTR_PT(282) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(284) OR ROM64_INSTR_PT(285)
     OR ROM64_INSTR_PT(287) OR ROM64_INSTR_PT(290)
     OR ROM64_INSTR_PT(293) OR ROM64_INSTR_PT(294)
     OR ROM64_INSTR_PT(297) OR ROM64_INSTR_PT(298)
     OR ROM64_INSTR_PT(299) OR ROM64_INSTR_PT(302)
     OR ROM64_INSTR_PT(305) OR ROM64_INSTR_PT(308)
     OR ROM64_INSTR_PT(311) OR ROM64_INSTR_PT(315)
     OR ROM64_INSTR_PT(319) OR ROM64_INSTR_PT(331)
     OR ROM64_INSTR_PT(339) OR ROM64_INSTR_PT(348)
     OR ROM64_INSTR_PT(353) OR ROM64_INSTR_PT(364)
     OR ROM64_INSTR_PT(372) OR ROM64_INSTR_PT(374)
     OR ROM64_INSTR_PT(375) OR ROM64_INSTR_PT(379)
     OR ROM64_INSTR_PT(381) OR ROM64_INSTR_PT(383)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(385)
     OR ROM64_INSTR_PT(391) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(395) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(404) OR ROM64_INSTR_PT(405)
     OR ROM64_INSTR_PT(410) OR ROM64_INSTR_PT(413)
     OR ROM64_INSTR_PT(414) OR ROM64_INSTR_PT(415)
     OR ROM64_INSTR_PT(418) OR ROM64_INSTR_PT(424)
     OR ROM64_INSTR_PT(425) OR ROM64_INSTR_PT(426)
     OR ROM64_INSTR_PT(428) OR ROM64_INSTR_PT(429)
     OR ROM64_INSTR_PT(430) OR ROM64_INSTR_PT(432)
     OR ROM64_INSTR_PT(435) OR ROM64_INSTR_PT(437)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(451) OR ROM64_INSTR_PT(453)
     OR ROM64_INSTR_PT(456) OR ROM64_INSTR_PT(457)
     OR ROM64_INSTR_PT(460) OR ROM64_INSTR_PT(467)
     OR ROM64_INSTR_PT(473) OR ROM64_INSTR_PT(475)
     OR ROM64_INSTR_PT(478) OR ROM64_INSTR_PT(481)
     OR ROM64_INSTR_PT(482) OR ROM64_INSTR_PT(484)
     OR ROM64_INSTR_PT(485) OR ROM64_INSTR_PT(488)
     OR ROM64_INSTR_PT(490) OR ROM64_INSTR_PT(493)
     OR ROM64_INSTR_PT(495) OR ROM64_INSTR_PT(496)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(505)
     OR ROM64_INSTR_PT(506) OR ROM64_INSTR_PT(507)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(511)
     OR ROM64_INSTR_PT(512) OR ROM64_INSTR_PT(517)
     OR ROM64_INSTR_PT(521) OR ROM64_INSTR_PT(522)
     OR ROM64_INSTR_PT(525) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(531) OR ROM64_INSTR_PT(534)
     OR ROM64_INSTR_PT(539) OR ROM64_INSTR_PT(546)
     OR ROM64_INSTR_PT(552) OR ROM64_INSTR_PT(553)
     OR ROM64_INSTR_PT(554) OR ROM64_INSTR_PT(555)
     OR ROM64_INSTR_PT(557) OR ROM64_INSTR_PT(558)
     OR ROM64_INSTR_PT(559) OR ROM64_INSTR_PT(563)
     OR ROM64_INSTR_PT(564) OR ROM64_INSTR_PT(568)
     OR ROM64_INSTR_PT(569) OR ROM64_INSTR_PT(577)
     OR ROM64_INSTR_PT(579) OR ROM64_INSTR_PT(580)
     OR ROM64_INSTR_PT(582) OR ROM64_INSTR_PT(583)
     OR ROM64_INSTR_PT(588) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(592) OR ROM64_INSTR_PT(595)
     OR ROM64_INSTR_PT(597) OR ROM64_INSTR_PT(600)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(608)
     OR ROM64_INSTR_PT(611) OR ROM64_INSTR_PT(615)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(619)
     OR ROM64_INSTR_PT(623) OR ROM64_INSTR_PT(627)
     OR ROM64_INSTR_PT(629) OR ROM64_INSTR_PT(632)
     OR ROM64_INSTR_PT(633) OR ROM64_INSTR_PT(636)
     OR ROM64_INSTR_PT(639) OR ROM64_INSTR_PT(642)
     OR ROM64_INSTR_PT(643) OR ROM64_INSTR_PT(644)
     OR ROM64_INSTR_PT(655) OR ROM64_INSTR_PT(660)
     OR ROM64_INSTR_PT(664) OR ROM64_INSTR_PT(666)
     OR ROM64_INSTR_PT(678) OR ROM64_INSTR_PT(702)
     OR ROM64_INSTR_PT(713) OR ROM64_INSTR_PT(722)
     OR ROM64_INSTR_PT(728) OR ROM64_INSTR_PT(735)
     OR ROM64_INSTR_PT(736) OR ROM64_INSTR_PT(738)
     OR ROM64_INSTR_PT(739) OR ROM64_INSTR_PT(744)
     OR ROM64_INSTR_PT(761) OR ROM64_INSTR_PT(769)
     OR ROM64_INSTR_PT(770) OR ROM64_INSTR_PT(776)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(811)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(824)
     OR ROM64_INSTR_PT(832) OR ROM64_INSTR_PT(855)
     OR ROM64_INSTR_PT(856) OR ROM64_INSTR_PT(864)
     OR ROM64_INSTR_PT(870));
MQQ920:TEMPLATE(29) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(7)
     OR ROM64_INSTR_PT(8) OR ROM64_INSTR_PT(9)
     OR ROM64_INSTR_PT(11) OR ROM64_INSTR_PT(14)
     OR ROM64_INSTR_PT(15) OR ROM64_INSTR_PT(17)
     OR ROM64_INSTR_PT(18) OR ROM64_INSTR_PT(22)
     OR ROM64_INSTR_PT(25) OR ROM64_INSTR_PT(28)
     OR ROM64_INSTR_PT(31) OR ROM64_INSTR_PT(38)
     OR ROM64_INSTR_PT(41) OR ROM64_INSTR_PT(49)
     OR ROM64_INSTR_PT(51) OR ROM64_INSTR_PT(52)
     OR ROM64_INSTR_PT(53) OR ROM64_INSTR_PT(61)
     OR ROM64_INSTR_PT(64) OR ROM64_INSTR_PT(70)
     OR ROM64_INSTR_PT(71) OR ROM64_INSTR_PT(75)
     OR ROM64_INSTR_PT(76) OR ROM64_INSTR_PT(83)
     OR ROM64_INSTR_PT(86) OR ROM64_INSTR_PT(90)
     OR ROM64_INSTR_PT(93) OR ROM64_INSTR_PT(97)
     OR ROM64_INSTR_PT(99) OR ROM64_INSTR_PT(100)
     OR ROM64_INSTR_PT(102) OR ROM64_INSTR_PT(105)
     OR ROM64_INSTR_PT(113) OR ROM64_INSTR_PT(115)
     OR ROM64_INSTR_PT(116) OR ROM64_INSTR_PT(117)
     OR ROM64_INSTR_PT(124) OR ROM64_INSTR_PT(127)
     OR ROM64_INSTR_PT(132) OR ROM64_INSTR_PT(133)
     OR ROM64_INSTR_PT(134) OR ROM64_INSTR_PT(136)
     OR ROM64_INSTR_PT(137) OR ROM64_INSTR_PT(140)
     OR ROM64_INSTR_PT(144) OR ROM64_INSTR_PT(148)
     OR ROM64_INSTR_PT(153) OR ROM64_INSTR_PT(158)
     OR ROM64_INSTR_PT(164) OR ROM64_INSTR_PT(168)
     OR ROM64_INSTR_PT(169) OR ROM64_INSTR_PT(171)
     OR ROM64_INSTR_PT(172) OR ROM64_INSTR_PT(181)
     OR ROM64_INSTR_PT(184) OR ROM64_INSTR_PT(185)
     OR ROM64_INSTR_PT(186) OR ROM64_INSTR_PT(194)
     OR ROM64_INSTR_PT(199) OR ROM64_INSTR_PT(202)
     OR ROM64_INSTR_PT(204) OR ROM64_INSTR_PT(211)
     OR ROM64_INSTR_PT(215) OR ROM64_INSTR_PT(217)
     OR ROM64_INSTR_PT(218) OR ROM64_INSTR_PT(219)
     OR ROM64_INSTR_PT(222) OR ROM64_INSTR_PT(226)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(238) OR ROM64_INSTR_PT(241)
     OR ROM64_INSTR_PT(245) OR ROM64_INSTR_PT(252)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(263) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(270)
     OR ROM64_INSTR_PT(271) OR ROM64_INSTR_PT(272)
     OR ROM64_INSTR_PT(273) OR ROM64_INSTR_PT(275)
     OR ROM64_INSTR_PT(276) OR ROM64_INSTR_PT(277)
     OR ROM64_INSTR_PT(282) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(285) OR ROM64_INSTR_PT(287)
     OR ROM64_INSTR_PT(293) OR ROM64_INSTR_PT(294)
     OR ROM64_INSTR_PT(297) OR ROM64_INSTR_PT(298)
     OR ROM64_INSTR_PT(299) OR ROM64_INSTR_PT(302)
     OR ROM64_INSTR_PT(305) OR ROM64_INSTR_PT(308)
     OR ROM64_INSTR_PT(311) OR ROM64_INSTR_PT(312)
     OR ROM64_INSTR_PT(315) OR ROM64_INSTR_PT(319)
     OR ROM64_INSTR_PT(324) OR ROM64_INSTR_PT(325)
     OR ROM64_INSTR_PT(331) OR ROM64_INSTR_PT(340)
     OR ROM64_INSTR_PT(361) OR ROM64_INSTR_PT(364)
     OR ROM64_INSTR_PT(374) OR ROM64_INSTR_PT(375)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(383)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(385)
     OR ROM64_INSTR_PT(388) OR ROM64_INSTR_PT(391)
     OR ROM64_INSTR_PT(394) OR ROM64_INSTR_PT(401)
     OR ROM64_INSTR_PT(403) OR ROM64_INSTR_PT(404)
     OR ROM64_INSTR_PT(406) OR ROM64_INSTR_PT(410)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(424) OR ROM64_INSTR_PT(428)
     OR ROM64_INSTR_PT(430) OR ROM64_INSTR_PT(432)
     OR ROM64_INSTR_PT(434) OR ROM64_INSTR_PT(437)
     OR ROM64_INSTR_PT(438) OR ROM64_INSTR_PT(439)
     OR ROM64_INSTR_PT(440) OR ROM64_INSTR_PT(441)
     OR ROM64_INSTR_PT(443) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(453)
     OR ROM64_INSTR_PT(454) OR ROM64_INSTR_PT(455)
     OR ROM64_INSTR_PT(468) OR ROM64_INSTR_PT(478)
     OR ROM64_INSTR_PT(481) OR ROM64_INSTR_PT(482)
     OR ROM64_INSTR_PT(484) OR ROM64_INSTR_PT(485)
     OR ROM64_INSTR_PT(493) OR ROM64_INSTR_PT(495)
     OR ROM64_INSTR_PT(496) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(505)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(510)
     OR ROM64_INSTR_PT(511) OR ROM64_INSTR_PT(512)
     OR ROM64_INSTR_PT(516) OR ROM64_INSTR_PT(519)
     OR ROM64_INSTR_PT(521) OR ROM64_INSTR_PT(522)
     OR ROM64_INSTR_PT(525) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(531) OR ROM64_INSTR_PT(532)
     OR ROM64_INSTR_PT(534) OR ROM64_INSTR_PT(535)
     OR ROM64_INSTR_PT(544) OR ROM64_INSTR_PT(545)
     OR ROM64_INSTR_PT(546) OR ROM64_INSTR_PT(549)
     OR ROM64_INSTR_PT(552) OR ROM64_INSTR_PT(555)
     OR ROM64_INSTR_PT(558) OR ROM64_INSTR_PT(559)
     OR ROM64_INSTR_PT(563) OR ROM64_INSTR_PT(564)
     OR ROM64_INSTR_PT(566) OR ROM64_INSTR_PT(569)
     OR ROM64_INSTR_PT(571) OR ROM64_INSTR_PT(575)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(580) OR ROM64_INSTR_PT(581)
     OR ROM64_INSTR_PT(582) OR ROM64_INSTR_PT(583)
     OR ROM64_INSTR_PT(586) OR ROM64_INSTR_PT(587)
     OR ROM64_INSTR_PT(588) OR ROM64_INSTR_PT(589)
     OR ROM64_INSTR_PT(591) OR ROM64_INSTR_PT(595)
     OR ROM64_INSTR_PT(600) OR ROM64_INSTR_PT(604)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(607)
     OR ROM64_INSTR_PT(608) OR ROM64_INSTR_PT(615)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(625)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(628)
     OR ROM64_INSTR_PT(629) OR ROM64_INSTR_PT(632)
     OR ROM64_INSTR_PT(633) OR ROM64_INSTR_PT(639)
     OR ROM64_INSTR_PT(642) OR ROM64_INSTR_PT(644)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(664)
     OR ROM64_INSTR_PT(666) OR ROM64_INSTR_PT(678)
     OR ROM64_INSTR_PT(681) OR ROM64_INSTR_PT(698)
     OR ROM64_INSTR_PT(702) OR ROM64_INSTR_PT(722)
     OR ROM64_INSTR_PT(728) OR ROM64_INSTR_PT(731)
     OR ROM64_INSTR_PT(735) OR ROM64_INSTR_PT(738)
     OR ROM64_INSTR_PT(744) OR ROM64_INSTR_PT(761)
     OR ROM64_INSTR_PT(769) OR ROM64_INSTR_PT(776)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(832)
     OR ROM64_INSTR_PT(846) OR ROM64_INSTR_PT(854)
     OR ROM64_INSTR_PT(856) OR ROM64_INSTR_PT(864)
     OR ROM64_INSTR_PT(870));
MQQ921:TEMPLATE(30) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(5)
     OR ROM64_INSTR_PT(7) OR ROM64_INSTR_PT(9)
     OR ROM64_INSTR_PT(10) OR ROM64_INSTR_PT(14)
     OR ROM64_INSTR_PT(17) OR ROM64_INSTR_PT(21)
     OR ROM64_INSTR_PT(22) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(38) OR ROM64_INSTR_PT(41)
     OR ROM64_INSTR_PT(45) OR ROM64_INSTR_PT(50)
     OR ROM64_INSTR_PT(51) OR ROM64_INSTR_PT(52)
     OR ROM64_INSTR_PT(55) OR ROM64_INSTR_PT(61)
     OR ROM64_INSTR_PT(64) OR ROM64_INSTR_PT(70)
     OR ROM64_INSTR_PT(71) OR ROM64_INSTR_PT(75)
     OR ROM64_INSTR_PT(76) OR ROM64_INSTR_PT(77)
     OR ROM64_INSTR_PT(78) OR ROM64_INSTR_PT(80)
     OR ROM64_INSTR_PT(83) OR ROM64_INSTR_PT(84)
     OR ROM64_INSTR_PT(86) OR ROM64_INSTR_PT(89)
     OR ROM64_INSTR_PT(90) OR ROM64_INSTR_PT(92)
     OR ROM64_INSTR_PT(96) OR ROM64_INSTR_PT(99)
     OR ROM64_INSTR_PT(100) OR ROM64_INSTR_PT(102)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(105)
     OR ROM64_INSTR_PT(106) OR ROM64_INSTR_PT(110)
     OR ROM64_INSTR_PT(113) OR ROM64_INSTR_PT(114)
     OR ROM64_INSTR_PT(115) OR ROM64_INSTR_PT(116)
     OR ROM64_INSTR_PT(117) OR ROM64_INSTR_PT(118)
     OR ROM64_INSTR_PT(121) OR ROM64_INSTR_PT(124)
     OR ROM64_INSTR_PT(127) OR ROM64_INSTR_PT(132)
     OR ROM64_INSTR_PT(136) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(143)
     OR ROM64_INSTR_PT(144) OR ROM64_INSTR_PT(148)
     OR ROM64_INSTR_PT(153) OR ROM64_INSTR_PT(169)
     OR ROM64_INSTR_PT(171) OR ROM64_INSTR_PT(175)
     OR ROM64_INSTR_PT(177) OR ROM64_INSTR_PT(180)
     OR ROM64_INSTR_PT(181) OR ROM64_INSTR_PT(183)
     OR ROM64_INSTR_PT(184) OR ROM64_INSTR_PT(185)
     OR ROM64_INSTR_PT(186) OR ROM64_INSTR_PT(188)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(199)
     OR ROM64_INSTR_PT(202) OR ROM64_INSTR_PT(204)
     OR ROM64_INSTR_PT(208) OR ROM64_INSTR_PT(213)
     OR ROM64_INSTR_PT(214) OR ROM64_INSTR_PT(215)
     OR ROM64_INSTR_PT(217) OR ROM64_INSTR_PT(218)
     OR ROM64_INSTR_PT(221) OR ROM64_INSTR_PT(222)
     OR ROM64_INSTR_PT(223) OR ROM64_INSTR_PT(226)
     OR ROM64_INSTR_PT(229) OR ROM64_INSTR_PT(230)
     OR ROM64_INSTR_PT(233) OR ROM64_INSTR_PT(238)
     OR ROM64_INSTR_PT(241) OR ROM64_INSTR_PT(252)
     OR ROM64_INSTR_PT(258) OR ROM64_INSTR_PT(260)
     OR ROM64_INSTR_PT(263) OR ROM64_INSTR_PT(264)
     OR ROM64_INSTR_PT(268) OR ROM64_INSTR_PT(270)
     OR ROM64_INSTR_PT(271) OR ROM64_INSTR_PT(274)
     OR ROM64_INSTR_PT(275) OR ROM64_INSTR_PT(276)
     OR ROM64_INSTR_PT(280) OR ROM64_INSTR_PT(282)
     OR ROM64_INSTR_PT(285) OR ROM64_INSTR_PT(286)
     OR ROM64_INSTR_PT(293) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(298) OR ROM64_INSTR_PT(299)
     OR ROM64_INSTR_PT(302) OR ROM64_INSTR_PT(305)
     OR ROM64_INSTR_PT(308) OR ROM64_INSTR_PT(315)
     OR ROM64_INSTR_PT(319) OR ROM64_INSTR_PT(322)
     OR ROM64_INSTR_PT(331) OR ROM64_INSTR_PT(339)
     OR ROM64_INSTR_PT(347) OR ROM64_INSTR_PT(349)
     OR ROM64_INSTR_PT(350) OR ROM64_INSTR_PT(358)
     OR ROM64_INSTR_PT(364) OR ROM64_INSTR_PT(367)
     OR ROM64_INSTR_PT(369) OR ROM64_INSTR_PT(371)
     OR ROM64_INSTR_PT(374) OR ROM64_INSTR_PT(375)
     OR ROM64_INSTR_PT(378) OR ROM64_INSTR_PT(379)
     OR ROM64_INSTR_PT(383) OR ROM64_INSTR_PT(385)
     OR ROM64_INSTR_PT(391) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(397) OR ROM64_INSTR_PT(403)
     OR ROM64_INSTR_PT(404) OR ROM64_INSTR_PT(410)
     OR ROM64_INSTR_PT(413) OR ROM64_INSTR_PT(414)
     OR ROM64_INSTR_PT(415) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(422) OR ROM64_INSTR_PT(424)
     OR ROM64_INSTR_PT(427) OR ROM64_INSTR_PT(430)
     OR ROM64_INSTR_PT(432) OR ROM64_INSTR_PT(434)
     OR ROM64_INSTR_PT(435) OR ROM64_INSTR_PT(437)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(445)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(453)
     OR ROM64_INSTR_PT(461) OR ROM64_INSTR_PT(463)
     OR ROM64_INSTR_PT(466) OR ROM64_INSTR_PT(478)
     OR ROM64_INSTR_PT(481) OR ROM64_INSTR_PT(482)
     OR ROM64_INSTR_PT(484) OR ROM64_INSTR_PT(485)
     OR ROM64_INSTR_PT(493) OR ROM64_INSTR_PT(495)
     OR ROM64_INSTR_PT(496) OR ROM64_INSTR_PT(503)
     OR ROM64_INSTR_PT(504) OR ROM64_INSTR_PT(505)
     OR ROM64_INSTR_PT(509) OR ROM64_INSTR_PT(510)
     OR ROM64_INSTR_PT(511) OR ROM64_INSTR_PT(512)
     OR ROM64_INSTR_PT(521) OR ROM64_INSTR_PT(522)
     OR ROM64_INSTR_PT(523) OR ROM64_INSTR_PT(525)
     OR ROM64_INSTR_PT(534) OR ROM64_INSTR_PT(540)
     OR ROM64_INSTR_PT(545) OR ROM64_INSTR_PT(546)
     OR ROM64_INSTR_PT(552) OR ROM64_INSTR_PT(555)
     OR ROM64_INSTR_PT(557) OR ROM64_INSTR_PT(558)
     OR ROM64_INSTR_PT(559) OR ROM64_INSTR_PT(563)
     OR ROM64_INSTR_PT(569) OR ROM64_INSTR_PT(571)
     OR ROM64_INSTR_PT(576) OR ROM64_INSTR_PT(579)
     OR ROM64_INSTR_PT(582) OR ROM64_INSTR_PT(583)
     OR ROM64_INSTR_PT(584) OR ROM64_INSTR_PT(588)
     OR ROM64_INSTR_PT(591) OR ROM64_INSTR_PT(592)
     OR ROM64_INSTR_PT(595) OR ROM64_INSTR_PT(596)
     OR ROM64_INSTR_PT(600) OR ROM64_INSTR_PT(606)
     OR ROM64_INSTR_PT(608) OR ROM64_INSTR_PT(609)
     OR ROM64_INSTR_PT(613) OR ROM64_INSTR_PT(615)
     OR ROM64_INSTR_PT(618) OR ROM64_INSTR_PT(619)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(629)
     OR ROM64_INSTR_PT(632) OR ROM64_INSTR_PT(633)
     OR ROM64_INSTR_PT(639) OR ROM64_INSTR_PT(642)
     OR ROM64_INSTR_PT(644) OR ROM64_INSTR_PT(666)
     OR ROM64_INSTR_PT(678) OR ROM64_INSTR_PT(685)
     OR ROM64_INSTR_PT(687) OR ROM64_INSTR_PT(691)
     OR ROM64_INSTR_PT(695) OR ROM64_INSTR_PT(716)
     OR ROM64_INSTR_PT(722) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(728)
     OR ROM64_INSTR_PT(731) OR ROM64_INSTR_PT(733)
     OR ROM64_INSTR_PT(735) OR ROM64_INSTR_PT(736)
     OR ROM64_INSTR_PT(738) OR ROM64_INSTR_PT(744)
     OR ROM64_INSTR_PT(761) OR ROM64_INSTR_PT(769)
     OR ROM64_INSTR_PT(770) OR ROM64_INSTR_PT(776)
     OR ROM64_INSTR_PT(834) OR ROM64_INSTR_PT(846)
     OR ROM64_INSTR_PT(856) OR ROM64_INSTR_PT(864)
     OR ROM64_INSTR_PT(870));
MQQ922:TEMPLATE(31) <= 
    (ROM64_INSTR_PT(33) OR ROM64_INSTR_PT(60)
     OR ROM64_INSTR_PT(79) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(103) OR ROM64_INSTR_PT(142)
     OR ROM64_INSTR_PT(147) OR ROM64_INSTR_PT(150)
     OR ROM64_INSTR_PT(160) OR ROM64_INSTR_PT(168)
     OR ROM64_INSTR_PT(176) OR ROM64_INSTR_PT(187)
     OR ROM64_INSTR_PT(207) OR ROM64_INSTR_PT(209)
     OR ROM64_INSTR_PT(219) OR ROM64_INSTR_PT(224)
     OR ROM64_INSTR_PT(228) OR ROM64_INSTR_PT(231)
     OR ROM64_INSTR_PT(247) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(281) OR ROM64_INSTR_PT(288)
     OR ROM64_INSTR_PT(296) OR ROM64_INSTR_PT(304)
     OR ROM64_INSTR_PT(309) OR ROM64_INSTR_PT(314)
     OR ROM64_INSTR_PT(327) OR ROM64_INSTR_PT(332)
     OR ROM64_INSTR_PT(341) OR ROM64_INSTR_PT(352)
     OR ROM64_INSTR_PT(361) OR ROM64_INSTR_PT(374)
     OR ROM64_INSTR_PT(401) OR ROM64_INSTR_PT(406)
     OR ROM64_INSTR_PT(464) OR ROM64_INSTR_PT(471)
     OR ROM64_INSTR_PT(491) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(632) OR ROM64_INSTR_PT(635)
     OR ROM64_INSTR_PT(641) OR ROM64_INSTR_PT(654)
     OR ROM64_INSTR_PT(675) OR ROM64_INSTR_PT(723)
     OR ROM64_INSTR_PT(724) OR ROM64_INSTR_PT(728)
     OR ROM64_INSTR_PT(733) OR ROM64_INSTR_PT(735)
     OR ROM64_INSTR_PT(738) OR ROM64_INSTR_PT(759)
     OR ROM64_INSTR_PT(766) OR ROM64_INSTR_PT(781)
     OR ROM64_INSTR_PT(794) OR ROM64_INSTR_PT(809)
    );
MQQ923:UCODE_END <= 
    (ROM64_INSTR_PT(198) OR ROM64_INSTR_PT(200)
     OR ROM64_INSTR_PT(212) OR ROM64_INSTR_PT(386)
     OR ROM64_INSTR_PT(443) OR ROM64_INSTR_PT(444)
     OR ROM64_INSTR_PT(452) OR ROM64_INSTR_PT(516)
     OR ROM64_INSTR_PT(518) OR ROM64_INSTR_PT(528)
     OR ROM64_INSTR_PT(542) OR ROM64_INSTR_PT(550)
     OR ROM64_INSTR_PT(556) OR ROM64_INSTR_PT(560)
     OR ROM64_INSTR_PT(567) OR ROM64_INSTR_PT(574)
     OR ROM64_INSTR_PT(577) OR ROM64_INSTR_PT(578)
     OR ROM64_INSTR_PT(581) OR ROM64_INSTR_PT(593)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(606)
     OR ROM64_INSTR_PT(607) OR ROM64_INSTR_PT(622)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(668)
     OR ROM64_INSTR_PT(690) OR ROM64_INSTR_PT(699)
     OR ROM64_INSTR_PT(704) OR ROM64_INSTR_PT(706)
     OR ROM64_INSTR_PT(714) OR ROM64_INSTR_PT(718)
     OR ROM64_INSTR_PT(741) OR ROM64_INSTR_PT(785)
     OR ROM64_INSTR_PT(790) OR ROM64_INSTR_PT(813)
     OR ROM64_INSTR_PT(823) OR ROM64_INSTR_PT(824)
     OR ROM64_INSTR_PT(826) OR ROM64_INSTR_PT(828)
     OR ROM64_INSTR_PT(841) OR ROM64_INSTR_PT(844)
     OR ROM64_INSTR_PT(845) OR ROM64_INSTR_PT(849)
     OR ROM64_INSTR_PT(854));
MQQ924:UCODE_END_EARLY <= 
    (ROM64_INSTR_PT(376) OR ROM64_INSTR_PT(390)
     OR ROM64_INSTR_PT(650) OR ROM64_INSTR_PT(676)
     OR ROM64_INSTR_PT(683) OR ROM64_INSTR_PT(689)
     OR ROM64_INSTR_PT(730) OR ROM64_INSTR_PT(742)
     OR ROM64_INSTR_PT(757) OR ROM64_INSTR_PT(760)
     OR ROM64_INSTR_PT(787) OR ROM64_INSTR_PT(788)
     OR ROM64_INSTR_PT(800) OR ROM64_INSTR_PT(802)
     OR ROM64_INSTR_PT(803) OR ROM64_INSTR_PT(807)
     OR ROM64_INSTR_PT(814) OR ROM64_INSTR_PT(818)
     OR ROM64_INSTR_PT(825) OR ROM64_INSTR_PT(830)
     OR ROM64_INSTR_PT(874));
MQQ925:LOOP_BEGIN <= 
    (ROM64_INSTR_PT(26) OR ROM64_INSTR_PT(55)
     OR ROM64_INSTR_PT(104) OR ROM64_INSTR_PT(124)
     OR ROM64_INSTR_PT(147) OR ROM64_INSTR_PT(210)
     OR ROM64_INSTR_PT(228) OR ROM64_INSTR_PT(231)
     OR ROM64_INSTR_PT(239) OR ROM64_INSTR_PT(246)
     OR ROM64_INSTR_PT(255) OR ROM64_INSTR_PT(306)
     OR ROM64_INSTR_PT(310) OR ROM64_INSTR_PT(316)
     OR ROM64_INSTR_PT(322) OR ROM64_INSTR_PT(349)
     OR ROM64_INSTR_PT(369) OR ROM64_INSTR_PT(379)
     OR ROM64_INSTR_PT(411) OR ROM64_INSTR_PT(412)
     OR ROM64_INSTR_PT(436) OR ROM64_INSTR_PT(450)
     OR ROM64_INSTR_PT(462) OR ROM64_INSTR_PT(487)
     OR ROM64_INSTR_PT(493) OR ROM64_INSTR_PT(496)
     OR ROM64_INSTR_PT(546) OR ROM64_INSTR_PT(559)
     OR ROM64_INSTR_PT(572) OR ROM64_INSTR_PT(590)
     OR ROM64_INSTR_PT(610));
MQQ926:LOOP_END <= 
    (ROM64_INSTR_PT(149) OR ROM64_INSTR_PT(156)
     OR ROM64_INSTR_PT(376) OR ROM64_INSTR_PT(469)
     OR ROM64_INSTR_PT(494) OR ROM64_INSTR_PT(502)
     OR ROM64_INSTR_PT(565) OR ROM64_INSTR_PT(638)
     OR ROM64_INSTR_PT(647) OR ROM64_INSTR_PT(656)
     OR ROM64_INSTR_PT(680) OR ROM64_INSTR_PT(701)
     OR ROM64_INSTR_PT(751) OR ROM64_INSTR_PT(775)
     OR ROM64_INSTR_PT(779) OR ROM64_INSTR_PT(789)
     OR ROM64_INSTR_PT(799) OR ROM64_INSTR_PT(807)
     OR ROM64_INSTR_PT(815) OR ROM64_INSTR_PT(816)
     OR ROM64_INSTR_PT(850) OR ROM64_INSTR_PT(862)
     OR ROM64_INSTR_PT(875));
MQQ927:COUNT_SRC(0) <= 
    (ROM64_INSTR_PT(72) OR ROM64_INSTR_PT(752)
     OR ROM64_INSTR_PT(768) OR ROM64_INSTR_PT(876)
     OR ROM64_INSTR_PT(881) OR ROM64_INSTR_PT(882)
     OR ROM64_INSTR_PT(887) OR ROM64_INSTR_PT(888)
     OR ROM64_INSTR_PT(889));
MQQ928:COUNT_SRC(1) <= 
    (ROM64_INSTR_PT(839) OR ROM64_INSTR_PT(879)
     OR ROM64_INSTR_PT(882) OR ROM64_INSTR_PT(884)
     OR ROM64_INSTR_PT(885) OR ROM64_INSTR_PT(888)
     OR ROM64_INSTR_PT(889));
MQQ929:COUNT_SRC(2) <= 
    (ROM64_INSTR_PT(686) OR ROM64_INSTR_PT(752)
     OR ROM64_INSTR_PT(768) OR ROM64_INSTR_PT(831)
     OR ROM64_INSTR_PT(839) OR ROM64_INSTR_PT(887)
     OR ROM64_INSTR_PT(888) OR ROM64_INSTR_PT(889)
    );
MQQ930:EXTRT <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(6)
     OR ROM64_INSTR_PT(19) OR ROM64_INSTR_PT(24)
     OR ROM64_INSTR_PT(27) OR ROM64_INSTR_PT(47)
     OR ROM64_INSTR_PT(48) OR ROM64_INSTR_PT(63)
     OR ROM64_INSTR_PT(69) OR ROM64_INSTR_PT(74)
     OR ROM64_INSTR_PT(91) OR ROM64_INSTR_PT(95)
     OR ROM64_INSTR_PT(98) OR ROM64_INSTR_PT(107)
     OR ROM64_INSTR_PT(120) OR ROM64_INSTR_PT(123)
     OR ROM64_INSTR_PT(130) OR ROM64_INSTR_PT(131)
     OR ROM64_INSTR_PT(133) OR ROM64_INSTR_PT(135)
     OR ROM64_INSTR_PT(138) OR ROM64_INSTR_PT(140)
     OR ROM64_INSTR_PT(141) OR ROM64_INSTR_PT(151)
     OR ROM64_INSTR_PT(152) OR ROM64_INSTR_PT(159)
     OR ROM64_INSTR_PT(163) OR ROM64_INSTR_PT(164)
     OR ROM64_INSTR_PT(167) OR ROM64_INSTR_PT(189)
     OR ROM64_INSTR_PT(192) OR ROM64_INSTR_PT(220)
     OR ROM64_INSTR_PT(227) OR ROM64_INSTR_PT(234)
     OR ROM64_INSTR_PT(235) OR ROM64_INSTR_PT(250)
     OR ROM64_INSTR_PT(253) OR ROM64_INSTR_PT(258)
     OR ROM64_INSTR_PT(266) OR ROM64_INSTR_PT(267)
     OR ROM64_INSTR_PT(279) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(300) OR ROM64_INSTR_PT(301)
     OR ROM64_INSTR_PT(303) OR ROM64_INSTR_PT(317)
     OR ROM64_INSTR_PT(318) OR ROM64_INSTR_PT(328)
     OR ROM64_INSTR_PT(330) OR ROM64_INSTR_PT(331)
     OR ROM64_INSTR_PT(335) OR ROM64_INSTR_PT(337)
     OR ROM64_INSTR_PT(338) OR ROM64_INSTR_PT(344)
     OR ROM64_INSTR_PT(355) OR ROM64_INSTR_PT(356)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(393)
     OR ROM64_INSTR_PT(394) OR ROM64_INSTR_PT(398)
     OR ROM64_INSTR_PT(418) OR ROM64_INSTR_PT(423)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(447)
     OR ROM64_INSTR_PT(449) OR ROM64_INSTR_PT(476)
     OR ROM64_INSTR_PT(486) OR ROM64_INSTR_PT(487)
     OR ROM64_INSTR_PT(496) OR ROM64_INSTR_PT(500)
     OR ROM64_INSTR_PT(501) OR ROM64_INSTR_PT(526)
     OR ROM64_INSTR_PT(547) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(594) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(624) OR ROM64_INSTR_PT(630)
     OR ROM64_INSTR_PT(631) OR ROM64_INSTR_PT(640)
     OR ROM64_INSTR_PT(651) OR ROM64_INSTR_PT(665)
     OR ROM64_INSTR_PT(670) OR ROM64_INSTR_PT(671)
     OR ROM64_INSTR_PT(672) OR ROM64_INSTR_PT(673)
     OR ROM64_INSTR_PT(674) OR ROM64_INSTR_PT(688)
     OR ROM64_INSTR_PT(696) OR ROM64_INSTR_PT(700)
     OR ROM64_INSTR_PT(707) OR ROM64_INSTR_PT(712)
     OR ROM64_INSTR_PT(727) OR ROM64_INSTR_PT(732)
     OR ROM64_INSTR_PT(737) OR ROM64_INSTR_PT(743)
     OR ROM64_INSTR_PT(744) OR ROM64_INSTR_PT(746)
     OR ROM64_INSTR_PT(747) OR ROM64_INSTR_PT(750)
     OR ROM64_INSTR_PT(755) OR ROM64_INSTR_PT(756)
     OR ROM64_INSTR_PT(763) OR ROM64_INSTR_PT(764)
     OR ROM64_INSTR_PT(767) OR ROM64_INSTR_PT(771)
     OR ROM64_INSTR_PT(774) OR ROM64_INSTR_PT(776)
     OR ROM64_INSTR_PT(777) OR ROM64_INSTR_PT(780)
     OR ROM64_INSTR_PT(782) OR ROM64_INSTR_PT(783)
     OR ROM64_INSTR_PT(784) OR ROM64_INSTR_PT(786)
     OR ROM64_INSTR_PT(793) OR ROM64_INSTR_PT(795)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(810)
     OR ROM64_INSTR_PT(812) OR ROM64_INSTR_PT(820)
     OR ROM64_INSTR_PT(821) OR ROM64_INSTR_PT(833)
     OR ROM64_INSTR_PT(835) OR ROM64_INSTR_PT(837)
     OR ROM64_INSTR_PT(838) OR ROM64_INSTR_PT(848)
     OR ROM64_INSTR_PT(857) OR ROM64_INSTR_PT(859)
     OR ROM64_INSTR_PT(860) OR ROM64_INSTR_PT(863)
     OR ROM64_INSTR_PT(864) OR ROM64_INSTR_PT(865)
     OR ROM64_INSTR_PT(866) OR ROM64_INSTR_PT(867)
     OR ROM64_INSTR_PT(868) OR ROM64_INSTR_PT(871)
     OR ROM64_INSTR_PT(877) OR ROM64_INSTR_PT(878)
     OR ROM64_INSTR_PT(880));
MQQ931:EXTS1 <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(19)
     OR ROM64_INSTR_PT(32) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(47) OR ROM64_INSTR_PT(74)
     OR ROM64_INSTR_PT(81) OR ROM64_INSTR_PT(91)
     OR ROM64_INSTR_PT(94) OR ROM64_INSTR_PT(100)
     OR ROM64_INSTR_PT(131) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(138) OR ROM64_INSTR_PT(159)
     OR ROM64_INSTR_PT(165) OR ROM64_INSTR_PT(167)
     OR ROM64_INSTR_PT(193) OR ROM64_INSTR_PT(211)
     OR ROM64_INSTR_PT(225) OR ROM64_INSTR_PT(227)
     OR ROM64_INSTR_PT(232) OR ROM64_INSTR_PT(235)
     OR ROM64_INSTR_PT(279) OR ROM64_INSTR_PT(289)
     OR ROM64_INSTR_PT(291) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(300) OR ROM64_INSTR_PT(301)
     OR ROM64_INSTR_PT(317) OR ROM64_INSTR_PT(318)
     OR ROM64_INSTR_PT(326) OR ROM64_INSTR_PT(328)
     OR ROM64_INSTR_PT(330) OR ROM64_INSTR_PT(331)
     OR ROM64_INSTR_PT(335) OR ROM64_INSTR_PT(337)
     OR ROM64_INSTR_PT(338) OR ROM64_INSTR_PT(344)
     OR ROM64_INSTR_PT(350) OR ROM64_INSTR_PT(358)
     OR ROM64_INSTR_PT(373) OR ROM64_INSTR_PT(379)
     OR ROM64_INSTR_PT(393) OR ROM64_INSTR_PT(398)
     OR ROM64_INSTR_PT(400) OR ROM64_INSTR_PT(421)
     OR ROM64_INSTR_PT(438) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(449) OR ROM64_INSTR_PT(465)
     OR ROM64_INSTR_PT(476) OR ROM64_INSTR_PT(479)
     OR ROM64_INSTR_PT(486) OR ROM64_INSTR_PT(500)
     OR ROM64_INSTR_PT(526) OR ROM64_INSTR_PT(543)
     OR ROM64_INSTR_PT(566) OR ROM64_INSTR_PT(577)
     OR ROM64_INSTR_PT(581) OR ROM64_INSTR_PT(593)
     OR ROM64_INSTR_PT(594) OR ROM64_INSTR_PT(604)
     OR ROM64_INSTR_PT(624) OR ROM64_INSTR_PT(630)
     OR ROM64_INSTR_PT(631) OR ROM64_INSTR_PT(652)
     OR ROM64_INSTR_PT(669) OR ROM64_INSTR_PT(671)
     OR ROM64_INSTR_PT(672) OR ROM64_INSTR_PT(673)
     OR ROM64_INSTR_PT(674) OR ROM64_INSTR_PT(688)
     OR ROM64_INSTR_PT(692) OR ROM64_INSTR_PT(694)
     OR ROM64_INSTR_PT(697) OR ROM64_INSTR_PT(700)
     OR ROM64_INSTR_PT(707) OR ROM64_INSTR_PT(708)
     OR ROM64_INSTR_PT(710) OR ROM64_INSTR_PT(712)
     OR ROM64_INSTR_PT(715) OR ROM64_INSTR_PT(720)
     OR ROM64_INSTR_PT(725) OR ROM64_INSTR_PT(732)
     OR ROM64_INSTR_PT(737) OR ROM64_INSTR_PT(741)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(746)
     OR ROM64_INSTR_PT(747) OR ROM64_INSTR_PT(749)
     OR ROM64_INSTR_PT(750) OR ROM64_INSTR_PT(755)
     OR ROM64_INSTR_PT(758) OR ROM64_INSTR_PT(762)
     OR ROM64_INSTR_PT(763) OR ROM64_INSTR_PT(764)
     OR ROM64_INSTR_PT(767) OR ROM64_INSTR_PT(771)
     OR ROM64_INSTR_PT(774) OR ROM64_INSTR_PT(777)
     OR ROM64_INSTR_PT(778) OR ROM64_INSTR_PT(780)
     OR ROM64_INSTR_PT(782) OR ROM64_INSTR_PT(783)
     OR ROM64_INSTR_PT(784) OR ROM64_INSTR_PT(786)
     OR ROM64_INSTR_PT(793) OR ROM64_INSTR_PT(795)
     OR ROM64_INSTR_PT(796) OR ROM64_INSTR_PT(806)
     OR ROM64_INSTR_PT(810) OR ROM64_INSTR_PT(812)
     OR ROM64_INSTR_PT(817) OR ROM64_INSTR_PT(820)
     OR ROM64_INSTR_PT(821) OR ROM64_INSTR_PT(823)
     OR ROM64_INSTR_PT(828) OR ROM64_INSTR_PT(835)
     OR ROM64_INSTR_PT(836) OR ROM64_INSTR_PT(837)
     OR ROM64_INSTR_PT(838) OR ROM64_INSTR_PT(842)
     OR ROM64_INSTR_PT(843) OR ROM64_INSTR_PT(844)
     OR ROM64_INSTR_PT(847) OR ROM64_INSTR_PT(848)
     OR ROM64_INSTR_PT(849) OR ROM64_INSTR_PT(851)
     OR ROM64_INSTR_PT(853) OR ROM64_INSTR_PT(859)
     OR ROM64_INSTR_PT(861) OR ROM64_INSTR_PT(865)
     OR ROM64_INSTR_PT(866) OR ROM64_INSTR_PT(867)
     OR ROM64_INSTR_PT(871) OR ROM64_INSTR_PT(877)
     OR ROM64_INSTR_PT(880));
MQQ932:EXTS2 <= 
    (ROM64_INSTR_PT(23) OR ROM64_INSTR_PT(27)
     OR ROM64_INSTR_PT(44) OR ROM64_INSTR_PT(47)
     OR ROM64_INSTR_PT(88) OR ROM64_INSTR_PT(91)
     OR ROM64_INSTR_PT(131) OR ROM64_INSTR_PT(138)
     OR ROM64_INSTR_PT(140) OR ROM64_INSTR_PT(152)
     OR ROM64_INSTR_PT(167) OR ROM64_INSTR_PT(178)
     OR ROM64_INSTR_PT(182) OR ROM64_INSTR_PT(189)
     OR ROM64_INSTR_PT(211) OR ROM64_INSTR_PT(298)
     OR ROM64_INSTR_PT(318) OR ROM64_INSTR_PT(330)
     OR ROM64_INSTR_PT(331) OR ROM64_INSTR_PT(335)
     OR ROM64_INSTR_PT(337) OR ROM64_INSTR_PT(344)
     OR ROM64_INSTR_PT(346) OR ROM64_INSTR_PT(350)
     OR ROM64_INSTR_PT(356) OR ROM64_INSTR_PT(358)
     OR ROM64_INSTR_PT(373) OR ROM64_INSTR_PT(380)
     OR ROM64_INSTR_PT(384) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(400) OR ROM64_INSTR_PT(418)
     OR ROM64_INSTR_PT(432) OR ROM64_INSTR_PT(441)
     OR ROM64_INSTR_PT(479) OR ROM64_INSTR_PT(500)
     OR ROM64_INSTR_PT(516) OR ROM64_INSTR_PT(526)
     OR ROM64_INSTR_PT(530) OR ROM64_INSTR_PT(542)
     OR ROM64_INSTR_PT(577) OR ROM64_INSTR_PT(580)
     OR ROM64_INSTR_PT(581) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(627)
     OR ROM64_INSTR_PT(631) OR ROM64_INSTR_PT(652)
     OR ROM64_INSTR_PT(672) OR ROM64_INSTR_PT(674)
     OR ROM64_INSTR_PT(696) OR ROM64_INSTR_PT(697)
     OR ROM64_INSTR_PT(700) OR ROM64_INSTR_PT(707)
     OR ROM64_INSTR_PT(715) OR ROM64_INSTR_PT(718)
     OR ROM64_INSTR_PT(725) OR ROM64_INSTR_PT(737)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(744)
     OR ROM64_INSTR_PT(745) OR ROM64_INSTR_PT(746)
     OR ROM64_INSTR_PT(750) OR ROM64_INSTR_PT(754)
     OR ROM64_INSTR_PT(756) OR ROM64_INSTR_PT(758)
     OR ROM64_INSTR_PT(763) OR ROM64_INSTR_PT(765)
     OR ROM64_INSTR_PT(767) OR ROM64_INSTR_PT(771)
     OR ROM64_INSTR_PT(772) OR ROM64_INSTR_PT(774)
     OR ROM64_INSTR_PT(776) OR ROM64_INSTR_PT(778)
     OR ROM64_INSTR_PT(784) OR ROM64_INSTR_PT(786)
     OR ROM64_INSTR_PT(812) OR ROM64_INSTR_PT(813)
     OR ROM64_INSTR_PT(820) OR ROM64_INSTR_PT(823)
     OR ROM64_INSTR_PT(828) OR ROM64_INSTR_PT(842)
     OR ROM64_INSTR_PT(843) OR ROM64_INSTR_PT(848)
     OR ROM64_INSTR_PT(854) OR ROM64_INSTR_PT(859)
     OR ROM64_INSTR_PT(860) OR ROM64_INSTR_PT(863)
     OR ROM64_INSTR_PT(866) OR ROM64_INSTR_PT(867)
     OR ROM64_INSTR_PT(868) OR ROM64_INSTR_PT(877)
     OR ROM64_INSTR_PT(880));
MQQ933:EXTS3 <= 
    (ROM64_INSTR_PT(47) OR ROM64_INSTR_PT(94)
     OR ROM64_INSTR_PT(100) OR ROM64_INSTR_PT(135)
     OR ROM64_INSTR_PT(159) OR ROM64_INSTR_PT(163)
     OR ROM64_INSTR_PT(192) OR ROM64_INSTR_PT(225)
     OR ROM64_INSTR_PT(235) OR ROM64_INSTR_PT(251)
     OR ROM64_INSTR_PT(279) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(300) OR ROM64_INSTR_PT(326)
     OR ROM64_INSTR_PT(337) OR ROM64_INSTR_PT(338)
     OR ROM64_INSTR_PT(350) OR ROM64_INSTR_PT(358)
     OR ROM64_INSTR_PT(379) OR ROM64_INSTR_PT(384)
     OR ROM64_INSTR_PT(398) OR ROM64_INSTR_PT(413)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(447)
     OR ROM64_INSTR_PT(524) OR ROM64_INSTR_PT(526)
     OR ROM64_INSTR_PT(561) OR ROM64_INSTR_PT(572)
     OR ROM64_INSTR_PT(594) OR ROM64_INSTR_PT(630)
     OR ROM64_INSTR_PT(670) OR ROM64_INSTR_PT(692)
     OR ROM64_INSTR_PT(697) OR ROM64_INSTR_PT(712)
     OR ROM64_INSTR_PT(715) OR ROM64_INSTR_PT(749)
     OR ROM64_INSTR_PT(758) OR ROM64_INSTR_PT(778)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(833)
     OR ROM64_INSTR_PT(837) OR ROM64_INSTR_PT(838)
     OR ROM64_INSTR_PT(871));
MQQ934:SEL0_5 <= 
    (ROM64_INSTR_PT(652) OR ROM64_INSTR_PT(718)
    );
MQQ935:SEL6_10(0) <= 
    (ROM64_INSTR_PT(40) OR ROM64_INSTR_PT(69)
     OR ROM64_INSTR_PT(82) OR ROM64_INSTR_PT(95)
     OR ROM64_INSTR_PT(107) OR ROM64_INSTR_PT(200)
     OR ROM64_INSTR_PT(211) OR ROM64_INSTR_PT(267)
     OR ROM64_INSTR_PT(386) OR ROM64_INSTR_PT(443)
     OR ROM64_INSTR_PT(444) OR ROM64_INSTR_PT(452)
     OR ROM64_INSTR_PT(516) OR ROM64_INSTR_PT(528)
     OR ROM64_INSTR_PT(529) OR ROM64_INSTR_PT(537)
     OR ROM64_INSTR_PT(542) OR ROM64_INSTR_PT(550)
     OR ROM64_INSTR_PT(560) OR ROM64_INSTR_PT(566)
     OR ROM64_INSTR_PT(573) OR ROM64_INSTR_PT(581)
     OR ROM64_INSTR_PT(604) OR ROM64_INSTR_PT(607)
     OR ROM64_INSTR_PT(621) OR ROM64_INSTR_PT(661)
     OR ROM64_INSTR_PT(698) OR ROM64_INSTR_PT(706)
     OR ROM64_INSTR_PT(790) OR ROM64_INSTR_PT(823)
     OR ROM64_INSTR_PT(854));
MQQ936:SEL6_10(1) <= 
    (ROM64_INSTR_PT(1) OR ROM64_INSTR_PT(3)
     OR ROM64_INSTR_PT(40) OR ROM64_INSTR_PT(54)
     OR ROM64_INSTR_PT(67) OR ROM64_INSTR_PT(69)
     OR ROM64_INSTR_PT(78) OR ROM64_INSTR_PT(82)
     OR ROM64_INSTR_PT(95) OR ROM64_INSTR_PT(107)
     OR ROM64_INSTR_PT(120) OR ROM64_INSTR_PT(182)
     OR ROM64_INSTR_PT(188) OR ROM64_INSTR_PT(256)
     OR ROM64_INSTR_PT(267) OR ROM64_INSTR_PT(287)
     OR ROM64_INSTR_PT(336) OR ROM64_INSTR_PT(346)
     OR ROM64_INSTR_PT(350) OR ROM64_INSTR_PT(354)
     OR ROM64_INSTR_PT(358) OR ROM64_INSTR_PT(380)
     OR ROM64_INSTR_PT(407) OR ROM64_INSTR_PT(431)
     OR ROM64_INSTR_PT(436) OR ROM64_INSTR_PT(459)
     OR ROM64_INSTR_PT(463) OR ROM64_INSTR_PT(487)
     OR ROM64_INSTR_PT(529) OR ROM64_INSTR_PT(530)
     OR ROM64_INSTR_PT(540) OR ROM64_INSTR_PT(580)
     OR ROM64_INSTR_PT(605) OR ROM64_INSTR_PT(640)
     OR ROM64_INSTR_PT(652) OR ROM64_INSTR_PT(658)
     OR ROM64_INSTR_PT(694) OR ROM64_INSTR_PT(697)
     OR ROM64_INSTR_PT(708) OR ROM64_INSTR_PT(715)
     OR ROM64_INSTR_PT(718) OR ROM64_INSTR_PT(720)
     OR ROM64_INSTR_PT(726) OR ROM64_INSTR_PT(727)
     OR ROM64_INSTR_PT(740) OR ROM64_INSTR_PT(769)
     OR ROM64_INSTR_PT(857) OR ROM64_INSTR_PT(864)
    );
MQQ937:SEL11_15(0) <= 
    (ROM64_INSTR_PT(37) OR ROM64_INSTR_PT(135)
     OR ROM64_INSTR_PT(193) OR ROM64_INSTR_PT(232)
     OR ROM64_INSTR_PT(248) OR ROM64_INSTR_PT(291)
     OR ROM64_INSTR_PT(373) OR ROM64_INSTR_PT(384)
     OR ROM64_INSTR_PT(438) OR ROM64_INSTR_PT(447)
     OR ROM64_INSTR_PT(465) OR ROM64_INSTR_PT(593)
     OR ROM64_INSTR_PT(663) OR ROM64_INSTR_PT(741)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(829)
    );
MQQ938:SEL11_15(1) <= 
    (ROM64_INSTR_PT(24) OR ROM64_INSTR_PT(27)
     OR ROM64_INSTR_PT(37) OR ROM64_INSTR_PT(44)
     OR ROM64_INSTR_PT(48) OR ROM64_INSTR_PT(59)
     OR ROM64_INSTR_PT(62) OR ROM64_INSTR_PT(63)
     OR ROM64_INSTR_PT(85) OR ROM64_INSTR_PT(98)
     OR ROM64_INSTR_PT(105) OR ROM64_INSTR_PT(115)
     OR ROM64_INSTR_PT(123) OR ROM64_INSTR_PT(130)
     OR ROM64_INSTR_PT(133) OR ROM64_INSTR_PT(140)
     OR ROM64_INSTR_PT(141) OR ROM64_INSTR_PT(151)
     OR ROM64_INSTR_PT(164) OR ROM64_INSTR_PT(189)
     OR ROM64_INSTR_PT(192) OR ROM64_INSTR_PT(193)
     OR ROM64_INSTR_PT(200) OR ROM64_INSTR_PT(220)
     OR ROM64_INSTR_PT(232) OR ROM64_INSTR_PT(234)
     OR ROM64_INSTR_PT(250) OR ROM64_INSTR_PT(253)
     OR ROM64_INSTR_PT(266) OR ROM64_INSTR_PT(283)
     OR ROM64_INSTR_PT(291) OR ROM64_INSTR_PT(303)
     OR ROM64_INSTR_PT(323) OR ROM64_INSTR_PT(354)
     OR ROM64_INSTR_PT(356) OR ROM64_INSTR_PT(373)
     OR ROM64_INSTR_PT(386) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(418) OR ROM64_INSTR_PT(423)
     OR ROM64_INSTR_PT(432) OR ROM64_INSTR_PT(438)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(444)
     OR ROM64_INSTR_PT(452) OR ROM64_INSTR_PT(465)
     OR ROM64_INSTR_PT(492) OR ROM64_INSTR_PT(516)
     OR ROM64_INSTR_PT(524) OR ROM64_INSTR_PT(528)
     OR ROM64_INSTR_PT(547) OR ROM64_INSTR_PT(550)
     OR ROM64_INSTR_PT(560) OR ROM64_INSTR_PT(573)
     OR ROM64_INSTR_PT(577) OR ROM64_INSTR_PT(591)
     OR ROM64_INSTR_PT(593) OR ROM64_INSTR_PT(597)
     OR ROM64_INSTR_PT(607) OR ROM64_INSTR_PT(621)
     OR ROM64_INSTR_PT(627) OR ROM64_INSTR_PT(634)
     OR ROM64_INSTR_PT(665) OR ROM64_INSTR_PT(698)
     OR ROM64_INSTR_PT(706) OR ROM64_INSTR_PT(717)
     OR ROM64_INSTR_PT(718) OR ROM64_INSTR_PT(734)
     OR ROM64_INSTR_PT(790) OR ROM64_INSTR_PT(806)
     OR ROM64_INSTR_PT(813) OR ROM64_INSTR_PT(824)
     OR ROM64_INSTR_PT(828) OR ROM64_INSTR_PT(840)
     OR ROM64_INSTR_PT(844) OR ROM64_INSTR_PT(849)
    );
MQQ939:SEL16_20(0) <= 
    (ROM64_INSTR_PT(6) OR ROM64_INSTR_PT(135)
     OR ROM64_INSTR_PT(194) OR ROM64_INSTR_PT(258)
     OR ROM64_INSTR_PT(260) OR ROM64_INSTR_PT(355)
     OR ROM64_INSTR_PT(447) OR ROM64_INSTR_PT(533)
     OR ROM64_INSTR_PT(798) OR ROM64_INSTR_PT(829)
    );
MQQ940:SEL16_20(1) <= 
    (ROM64_INSTR_PT(4) OR ROM64_INSTR_PT(12)
     OR ROM64_INSTR_PT(16) OR ROM64_INSTR_PT(40)
     OR ROM64_INSTR_PT(46) OR ROM64_INSTR_PT(48)
     OR ROM64_INSTR_PT(69) OR ROM64_INSTR_PT(74)
     OR ROM64_INSTR_PT(82) OR ROM64_INSTR_PT(87)
     OR ROM64_INSTR_PT(95) OR ROM64_INSTR_PT(100)
     OR ROM64_INSTR_PT(107) OR ROM64_INSTR_PT(126)
     OR ROM64_INSTR_PT(133) OR ROM64_INSTR_PT(135)
     OR ROM64_INSTR_PT(137) OR ROM64_INSTR_PT(141)
     OR ROM64_INSTR_PT(159) OR ROM64_INSTR_PT(164)
     OR ROM64_INSTR_PT(200) OR ROM64_INSTR_PT(204)
     OR ROM64_INSTR_PT(225) OR ROM64_INSTR_PT(251)
     OR ROM64_INSTR_PT(266) OR ROM64_INSTR_PT(267)
     OR ROM64_INSTR_PT(279) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(300) OR ROM64_INSTR_PT(319)
     OR ROM64_INSTR_PT(321) OR ROM64_INSTR_PT(336)
     OR ROM64_INSTR_PT(354) OR ROM64_INSTR_PT(355)
     OR ROM64_INSTR_PT(362) OR ROM64_INSTR_PT(379)
     OR ROM64_INSTR_PT(398) OR ROM64_INSTR_PT(413)
     OR ROM64_INSTR_PT(423) OR ROM64_INSTR_PT(444)
     OR ROM64_INSTR_PT(446) OR ROM64_INSTR_PT(447)
     OR ROM64_INSTR_PT(452) OR ROM64_INSTR_PT(470)
     OR ROM64_INSTR_PT(496) OR ROM64_INSTR_PT(513)
     OR ROM64_INSTR_PT(524) OR ROM64_INSTR_PT(528)
     OR ROM64_INSTR_PT(529) OR ROM64_INSTR_PT(541)
     OR ROM64_INSTR_PT(550) OR ROM64_INSTR_PT(560)
     OR ROM64_INSTR_PT(561) OR ROM64_INSTR_PT(566)
     OR ROM64_INSTR_PT(572) OR ROM64_INSTR_PT(573)
     OR ROM64_INSTR_PT(606) OR ROM64_INSTR_PT(607)
     OR ROM64_INSTR_PT(615) OR ROM64_INSTR_PT(621)
     OR ROM64_INSTR_PT(634) OR ROM64_INSTR_PT(648)
     OR ROM64_INSTR_PT(661) OR ROM64_INSTR_PT(698)
     OR ROM64_INSTR_PT(706) OR ROM64_INSTR_PT(717)
     OR ROM64_INSTR_PT(729) OR ROM64_INSTR_PT(773)
     OR ROM64_INSTR_PT(790) OR ROM64_INSTR_PT(798)
     OR ROM64_INSTR_PT(829) OR ROM64_INSTR_PT(838)
    );
MQQ941:SEL21_25(0) <= 
    (ROM64_INSTR_PT(197));
MQQ942:SEL21_25(1) <= 
    (ROM64_INSTR_PT(16) OR ROM64_INSTR_PT(46)
     OR ROM64_INSTR_PT(48) OR ROM64_INSTR_PT(63)
     OR ROM64_INSTR_PT(74) OR ROM64_INSTR_PT(87)
     OR ROM64_INSTR_PT(141) OR ROM64_INSTR_PT(200)
     OR ROM64_INSTR_PT(225) OR ROM64_INSTR_PT(266)
     OR ROM64_INSTR_PT(321) OR ROM64_INSTR_PT(354)
     OR ROM64_INSTR_PT(362) OR ROM64_INSTR_PT(423)
     OR ROM64_INSTR_PT(452) OR ROM64_INSTR_PT(470)
     OR ROM64_INSTR_PT(515) OR ROM64_INSTR_PT(528)
     OR ROM64_INSTR_PT(541) OR ROM64_INSTR_PT(550)
     OR ROM64_INSTR_PT(560) OR ROM64_INSTR_PT(572)
     OR ROM64_INSTR_PT(573) OR ROM64_INSTR_PT(634)
     OR ROM64_INSTR_PT(652) OR ROM64_INSTR_PT(706)
     OR ROM64_INSTR_PT(718) OR ROM64_INSTR_PT(729)
     OR ROM64_INSTR_PT(734) OR ROM64_INSTR_PT(790)
    );
MQQ943:SEL26_30 <= 
    (ROM64_INSTR_PT(16) OR ROM64_INSTR_PT(46)
     OR ROM64_INSTR_PT(48) OR ROM64_INSTR_PT(63)
     OR ROM64_INSTR_PT(74) OR ROM64_INSTR_PT(87)
     OR ROM64_INSTR_PT(141) OR ROM64_INSTR_PT(200)
     OR ROM64_INSTR_PT(225) OR ROM64_INSTR_PT(266)
     OR ROM64_INSTR_PT(321) OR ROM64_INSTR_PT(354)
     OR ROM64_INSTR_PT(362) OR ROM64_INSTR_PT(423)
     OR ROM64_INSTR_PT(452) OR ROM64_INSTR_PT(470)
     OR ROM64_INSTR_PT(515) OR ROM64_INSTR_PT(528)
     OR ROM64_INSTR_PT(541) OR ROM64_INSTR_PT(550)
     OR ROM64_INSTR_PT(560) OR ROM64_INSTR_PT(572)
     OR ROM64_INSTR_PT(573) OR ROM64_INSTR_PT(634)
     OR ROM64_INSTR_PT(652) OR ROM64_INSTR_PT(706)
     OR ROM64_INSTR_PT(718) OR ROM64_INSTR_PT(729)
     OR ROM64_INSTR_PT(734) OR ROM64_INSTR_PT(790)
    );
MQQ944:SEL31 <= 
    (ROM64_INSTR_PT(16) OR ROM64_INSTR_PT(46)
     OR ROM64_INSTR_PT(63) OR ROM64_INSTR_PT(74)
     OR ROM64_INSTR_PT(87) OR ROM64_INSTR_PT(141)
     OR ROM64_INSTR_PT(200) OR ROM64_INSTR_PT(266)
     OR ROM64_INSTR_PT(321) OR ROM64_INSTR_PT(350)
     OR ROM64_INSTR_PT(354) OR ROM64_INSTR_PT(358)
     OR ROM64_INSTR_PT(362) OR ROM64_INSTR_PT(423)
     OR ROM64_INSTR_PT(452) OR ROM64_INSTR_PT(470)
     OR ROM64_INSTR_PT(541) OR ROM64_INSTR_PT(542)
     OR ROM64_INSTR_PT(560) OR ROM64_INSTR_PT(561)
     OR ROM64_INSTR_PT(573) OR ROM64_INSTR_PT(634)
     OR ROM64_INSTR_PT(652) OR ROM64_INSTR_PT(697)
     OR ROM64_INSTR_PT(706) OR ROM64_INSTR_PT(715)
     OR ROM64_INSTR_PT(718) OR ROM64_INSTR_PT(729)
     OR ROM64_INSTR_PT(790) OR ROM64_INSTR_PT(823)
    );
MQQ945:CR_BF2FXM <= 
    (ROM64_INSTR_PT(717));
MQQ946:SKIP_COND <= 
    (ROM64_INSTR_PT(23) OR ROM64_INSTR_PT(34)
     OR ROM64_INSTR_PT(81) OR ROM64_INSTR_PT(88)
     OR ROM64_INSTR_PT(91) OR ROM64_INSTR_PT(127)
     OR ROM64_INSTR_PT(298) OR ROM64_INSTR_PT(330)
     OR ROM64_INSTR_PT(331) OR ROM64_INSTR_PT(335)
     OR ROM64_INSTR_PT(344) OR ROM64_INSTR_PT(369)
     OR ROM64_INSTR_PT(489) OR ROM64_INSTR_PT(662)
     OR ROM64_INSTR_PT(667) OR ROM64_INSTR_PT(677)
     OR ROM64_INSTR_PT(684) OR ROM64_INSTR_PT(725)
     OR ROM64_INSTR_PT(744) OR ROM64_INSTR_PT(745)
     OR ROM64_INSTR_PT(746) OR ROM64_INSTR_PT(747)
     OR ROM64_INSTR_PT(748) OR ROM64_INSTR_PT(750)
     OR ROM64_INSTR_PT(754) OR ROM64_INSTR_PT(755)
     OR ROM64_INSTR_PT(756) OR ROM64_INSTR_PT(765)
     OR ROM64_INSTR_PT(776) OR ROM64_INSTR_PT(782)
     OR ROM64_INSTR_PT(783) OR ROM64_INSTR_PT(784)
     OR ROM64_INSTR_PT(792) OR ROM64_INSTR_PT(795)
     OR ROM64_INSTR_PT(796) OR ROM64_INSTR_PT(804)
     OR ROM64_INSTR_PT(817) OR ROM64_INSTR_PT(819)
     OR ROM64_INSTR_PT(820) OR ROM64_INSTR_PT(821)
     OR ROM64_INSTR_PT(827) OR ROM64_INSTR_PT(842)
     OR ROM64_INSTR_PT(859) OR ROM64_INSTR_PT(867)
    );
MQQ947:SKIP_ZERO <= 
    (ROM64_INSTR_PT(301) OR ROM64_INSTR_PT(319)
     OR ROM64_INSTR_PT(393) OR ROM64_INSTR_PT(436)
     OR ROM64_INSTR_PT(487) OR ROM64_INSTR_PT(496)
     OR ROM64_INSTR_PT(778));
MQQ948:LOOP_ADDR(0) <= 
    (ROM64_INSTR_PT(235) OR ROM64_INSTR_PT(289)
     OR ROM64_INSTR_PT(301) OR ROM64_INSTR_PT(317)
     OR ROM64_INSTR_PT(328) OR ROM64_INSTR_PT(373)
     OR ROM64_INSTR_PT(479) OR ROM64_INSTR_PT(526)
     OR ROM64_INSTR_PT(674) OR ROM64_INSTR_PT(692)
     OR ROM64_INSTR_PT(700) OR ROM64_INSTR_PT(732)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(777)
     OR ROM64_INSTR_PT(778) OR ROM64_INSTR_PT(784)
     OR ROM64_INSTR_PT(837) OR ROM64_INSTR_PT(861)
     OR ROM64_INSTR_PT(866) OR ROM64_INSTR_PT(867)
    );
MQQ949:LOOP_ADDR(1) <= 
    (ROM64_INSTR_PT(289) OR ROM64_INSTR_PT(479)
     OR ROM64_INSTR_PT(526) OR ROM64_INSTR_PT(674)
     OR ROM64_INSTR_PT(732) OR ROM64_INSTR_PT(777)
     OR ROM64_INSTR_PT(784) OR ROM64_INSTR_PT(833)
     OR ROM64_INSTR_PT(837) OR ROM64_INSTR_PT(859)
     OR ROM64_INSTR_PT(867));
MQQ950:LOOP_ADDR(2) <= 
    (ROM64_INSTR_PT(393) OR ROM64_INSTR_PT(449)
     OR ROM64_INSTR_PT(486) OR ROM64_INSTR_PT(700)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(748)
     OR ROM64_INSTR_PT(754) OR ROM64_INSTR_PT(764)
    );
MQQ951:LOOP_ADDR(3) <= 
    (ROM64_INSTR_PT(317) OR ROM64_INSTR_PT(328)
     OR ROM64_INSTR_PT(501) OR ROM64_INSTR_PT(672)
     OR ROM64_INSTR_PT(688) OR ROM64_INSTR_PT(700)
     OR ROM64_INSTR_PT(707) OR ROM64_INSTR_PT(725)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(765)
     OR ROM64_INSTR_PT(767) OR ROM64_INSTR_PT(777)
     OR ROM64_INSTR_PT(836) OR ROM64_INSTR_PT(837)
     OR ROM64_INSTR_PT(859) OR ROM64_INSTR_PT(867)
     OR ROM64_INSTR_PT(878));
MQQ952:LOOP_ADDR(4) <= 
    (ROM64_INSTR_PT(37) OR ROM64_INSTR_PT(289)
     OR ROM64_INSTR_PT(301) OR ROM64_INSTR_PT(328)
     OR ROM64_INSTR_PT(373) OR ROM64_INSTR_PT(400)
     OR ROM64_INSTR_PT(421) OR ROM64_INSTR_PT(449)
     OR ROM64_INSTR_PT(479) OR ROM64_INSTR_PT(700)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(748)
     OR ROM64_INSTR_PT(750) OR ROM64_INSTR_PT(754)
     OR ROM64_INSTR_PT(762) OR ROM64_INSTR_PT(784)
     OR ROM64_INSTR_PT(837) OR ROM64_INSTR_PT(866)
     OR ROM64_INSTR_PT(867));
MQQ953:LOOP_ADDR(5) <= 
    (ROM64_INSTR_PT(37) OR ROM64_INSTR_PT(235)
     OR ROM64_INSTR_PT(289) OR ROM64_INSTR_PT(421)
     OR ROM64_INSTR_PT(449) OR ROM64_INSTR_PT(526)
     OR ROM64_INSTR_PT(688) OR ROM64_INSTR_PT(725)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(764)
     OR ROM64_INSTR_PT(772) OR ROM64_INSTR_PT(861)
     OR ROM64_INSTR_PT(866));
MQQ954:LOOP_ADDR(6) <= 
    (ROM64_INSTR_PT(37) OR ROM64_INSTR_PT(163)
     OR ROM64_INSTR_PT(289) OR ROM64_INSTR_PT(317)
     OR ROM64_INSTR_PT(373) OR ROM64_INSTR_PT(486)
     OR ROM64_INSTR_PT(672) OR ROM64_INSTR_PT(696)
     OR ROM64_INSTR_PT(700) OR ROM64_INSTR_PT(748)
     OR ROM64_INSTR_PT(750) OR ROM64_INSTR_PT(764)
     OR ROM64_INSTR_PT(767) OR ROM64_INSTR_PT(833)
     OR ROM64_INSTR_PT(837) OR ROM64_INSTR_PT(859)
     OR ROM64_INSTR_PT(861) OR ROM64_INSTR_PT(868)
    );
MQQ955:LOOP_ADDR(7) <= 
    (ROM64_INSTR_PT(37) OR ROM64_INSTR_PT(289)
     OR ROM64_INSTR_PT(301) OR ROM64_INSTR_PT(317)
     OR ROM64_INSTR_PT(328) OR ROM64_INSTR_PT(400)
     OR ROM64_INSTR_PT(421) OR ROM64_INSTR_PT(486)
     OR ROM64_INSTR_PT(651) OR ROM64_INSTR_PT(672)
     OR ROM64_INSTR_PT(674) OR ROM64_INSTR_PT(692)
     OR ROM64_INSTR_PT(725) OR ROM64_INSTR_PT(732)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(748)
     OR ROM64_INSTR_PT(777) OR ROM64_INSTR_PT(861)
     OR ROM64_INSTR_PT(867));
MQQ956:LOOP_ADDR(8) <= 
    (ROM64_INSTR_PT(400) OR ROM64_INSTR_PT(421)
     OR ROM64_INSTR_PT(449) OR ROM64_INSTR_PT(479)
     OR ROM64_INSTR_PT(486) OR ROM64_INSTR_PT(672)
     OR ROM64_INSTR_PT(696) OR ROM64_INSTR_PT(700)
     OR ROM64_INSTR_PT(707) OR ROM64_INSTR_PT(725)
     OR ROM64_INSTR_PT(748) OR ROM64_INSTR_PT(750)
     OR ROM64_INSTR_PT(754) OR ROM64_INSTR_PT(762)
     OR ROM64_INSTR_PT(764) OR ROM64_INSTR_PT(777)
     OR ROM64_INSTR_PT(861) OR ROM64_INSTR_PT(866)
    );
MQQ957:LOOP_ADDR(9) <= 
    (ROM64_INSTR_PT(301) OR ROM64_INSTR_PT(317)
     OR ROM64_INSTR_PT(328) OR ROM64_INSTR_PT(373)
     OR ROM64_INSTR_PT(393) OR ROM64_INSTR_PT(449)
     OR ROM64_INSTR_PT(486) OR ROM64_INSTR_PT(692)
     OR ROM64_INSTR_PT(743) OR ROM64_INSTR_PT(764)
     OR ROM64_INSTR_PT(772) OR ROM64_INSTR_PT(778)
     OR ROM64_INSTR_PT(784) OR ROM64_INSTR_PT(836)
     OR ROM64_INSTR_PT(837) OR ROM64_INSTR_PT(861)
    );
MQQ958:LOOP_INIT(0) <= 
    (ROM64_INSTR_PT(235) OR ROM64_INSTR_PT(369)
     OR ROM64_INSTR_PT(398) OR ROM64_INSTR_PT(572)
     OR ROM64_INSTR_PT(673) OR ROM64_INSTR_PT(692)
     OR ROM64_INSTR_PT(783) OR ROM64_INSTR_PT(795)
     OR ROM64_INSTR_PT(810) OR ROM64_INSTR_PT(817)
     OR ROM64_INSTR_PT(821) OR ROM64_INSTR_PT(837)
     OR ROM64_INSTR_PT(859) OR ROM64_INSTR_PT(867)
    );
MQQ959:LOOP_INIT(1) <= 
    (ROM64_INSTR_PT(890));
MQQ960:LOOP_INIT(2) <= 
    (ROM64_INSTR_PT(783) OR ROM64_INSTR_PT(817)
     OR ROM64_INSTR_PT(859) OR ROM64_INSTR_PT(867)
    );
MQQ961:EP <= 
    (ROM64_INSTR_PT(44) OR ROM64_INSTR_PT(59)
     OR ROM64_INSTR_PT(115) OR ROM64_INSTR_PT(137)
     OR ROM64_INSTR_PT(279) OR ROM64_INSTR_PT(297)
     OR ROM64_INSTR_PT(356) OR ROM64_INSTR_PT(394)
     OR ROM64_INSTR_PT(398) OR ROM64_INSTR_PT(432)
     OR ROM64_INSTR_PT(441) OR ROM64_INSTR_PT(446)
     OR ROM64_INSTR_PT(524) OR ROM64_INSTR_PT(561)
    );

end generate;
c32: if (regmode = 5) generate
begin

ROM64_INSTR_PT  <=  (others => '0');
rom_unused  <=  or_reduce(ROM64_INSTR_PT);
MQQ962:ROM32_INSTR_PT(1) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100000000"));
MQQ963:ROM32_INSTR_PT(2) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000000"));
MQQ964:ROM32_INSTR_PT(3) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000000"));
MQQ965:ROM32_INSTR_PT(4) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000000"));
MQQ966:ROM32_INSTR_PT(5) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110000000"));
MQQ967:ROM32_INSTR_PT(6) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000000"));
MQQ968:ROM32_INSTR_PT(7) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00100000"));
MQQ969:ROM32_INSTR_PT(8) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100000"));
MQQ970:ROM32_INSTR_PT(9) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100000"));
MQQ971:ROM32_INSTR_PT(10) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100000"));
MQQ972:ROM32_INSTR_PT(11) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000000"));
MQQ973:ROM32_INSTR_PT(12) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000000"));
MQQ974:ROM32_INSTR_PT(13) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010000"));
MQQ975:ROM32_INSTR_PT(14) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010000"));
MQQ976:ROM32_INSTR_PT(15) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101010000"));
MQQ977:ROM32_INSTR_PT(16) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110000"));
MQQ978:ROM32_INSTR_PT(17) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110000"));
MQQ979:ROM32_INSTR_PT(18) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011110000"));
MQQ980:ROM32_INSTR_PT(19) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110000"));
MQQ981:ROM32_INSTR_PT(20) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ982:ROM32_INSTR_PT(21) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010000"));
MQQ983:ROM32_INSTR_PT(22) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110000"));
MQQ984:ROM32_INSTR_PT(23) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ985:ROM32_INSTR_PT(24) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000000"));
MQQ986:ROM32_INSTR_PT(25) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100000"));
MQQ987:ROM32_INSTR_PT(26) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010000"));
MQQ988:ROM32_INSTR_PT(27) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010000"));
MQQ989:ROM32_INSTR_PT(28) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110000"));
MQQ990:ROM32_INSTR_PT(29) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ991:ROM32_INSTR_PT(30) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110000"));
MQQ992:ROM32_INSTR_PT(31) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010000"));
MQQ993:ROM32_INSTR_PT(32) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010000"));
MQQ994:ROM32_INSTR_PT(33) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110000"));
MQQ995:ROM32_INSTR_PT(34) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001000"));
MQQ996:ROM32_INSTR_PT(35) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001000"));
MQQ997:ROM32_INSTR_PT(36) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101001000"));
MQQ998:ROM32_INSTR_PT(37) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110001000"));
MQQ999:ROM32_INSTR_PT(38) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001000"));
MQQ1000:ROM32_INSTR_PT(39) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100101000"));
MQQ1001:ROM32_INSTR_PT(40) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101000"));
MQQ1002:ROM32_INSTR_PT(41) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001101000"));
MQQ1003:ROM32_INSTR_PT(42) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101000"));
MQQ1004:ROM32_INSTR_PT(43) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101000"));
MQQ1005:ROM32_INSTR_PT(44) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101000"));
MQQ1006:ROM32_INSTR_PT(45) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111101000"));
MQQ1007:ROM32_INSTR_PT(46) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001000"));
MQQ1008:ROM32_INSTR_PT(47) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101000"));
MQQ1009:ROM32_INSTR_PT(48) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001011000"));
MQQ1010:ROM32_INSTR_PT(49) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011011000"));
MQQ1011:ROM32_INSTR_PT(50) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011011000"));
MQQ1012:ROM32_INSTR_PT(51) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111000"));
MQQ1013:ROM32_INSTR_PT(52) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111000"));
MQQ1014:ROM32_INSTR_PT(53) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111000"));
MQQ1015:ROM32_INSTR_PT(54) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010011000"));
MQQ1016:ROM32_INSTR_PT(55) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111000"));
MQQ1017:ROM32_INSTR_PT(56) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111000"));
MQQ1018:ROM32_INSTR_PT(57) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111000"));
MQQ1019:ROM32_INSTR_PT(58) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111000"));
MQQ1020:ROM32_INSTR_PT(59) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001000"));
MQQ1021:ROM32_INSTR_PT(60) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001000"));
MQQ1022:ROM32_INSTR_PT(61) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011000"));
MQQ1023:ROM32_INSTR_PT(62) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011000"));
MQQ1024:ROM32_INSTR_PT(63) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100111000"));
MQQ1025:ROM32_INSTR_PT(64) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111000"));
MQQ1026:ROM32_INSTR_PT(65) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000000"));
MQQ1027:ROM32_INSTR_PT(66) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000000"));
MQQ1028:ROM32_INSTR_PT(67) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000000"));
MQQ1029:ROM32_INSTR_PT(68) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000000"));
MQQ1030:ROM32_INSTR_PT(69) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010000"));
MQQ1031:ROM32_INSTR_PT(70) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010000"));
MQQ1032:ROM32_INSTR_PT(71) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ1033:ROM32_INSTR_PT(72) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010000"));
MQQ1034:ROM32_INSTR_PT(73) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001000"));
MQQ1035:ROM32_INSTR_PT(74) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011000"));
MQQ1036:ROM32_INSTR_PT(75) <=
    Eq(( ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000"));
MQQ1037:ROM32_INSTR_PT(76) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000100"));
MQQ1038:ROM32_INSTR_PT(77) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000100"));
MQQ1039:ROM32_INSTR_PT(78) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000100"));
MQQ1040:ROM32_INSTR_PT(79) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000100"));
MQQ1041:ROM32_INSTR_PT(80) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000100"));
MQQ1042:ROM32_INSTR_PT(81) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000100"));
MQQ1043:ROM32_INSTR_PT(82) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100100"));
MQQ1044:ROM32_INSTR_PT(83) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100100"));
MQQ1045:ROM32_INSTR_PT(84) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100100"));
MQQ1046:ROM32_INSTR_PT(85) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11100100"));
MQQ1047:ROM32_INSTR_PT(86) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100100"));
MQQ1048:ROM32_INSTR_PT(87) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000100"));
MQQ1049:ROM32_INSTR_PT(88) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10000100"));
MQQ1050:ROM32_INSTR_PT(89) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100100"));
MQQ1051:ROM32_INSTR_PT(90) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110010100"));
MQQ1052:ROM32_INSTR_PT(91) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010100"));
MQQ1053:ROM32_INSTR_PT(92) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010100"));
MQQ1054:ROM32_INSTR_PT(93) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010100"));
MQQ1055:ROM32_INSTR_PT(94) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110100"));
MQQ1056:ROM32_INSTR_PT(95) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110100"));
MQQ1057:ROM32_INSTR_PT(96) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110100"));
MQQ1058:ROM32_INSTR_PT(97) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110100"));
MQQ1059:ROM32_INSTR_PT(98) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010100"));
MQQ1060:ROM32_INSTR_PT(99) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110100"));
MQQ1061:ROM32_INSTR_PT(100) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110100"));
MQQ1062:ROM32_INSTR_PT(101) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110100"));
MQQ1063:ROM32_INSTR_PT(102) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000100"));
MQQ1064:ROM32_INSTR_PT(103) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000100"));
MQQ1065:ROM32_INSTR_PT(104) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010100"));
MQQ1066:ROM32_INSTR_PT(105) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110100"));
MQQ1067:ROM32_INSTR_PT(106) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010100"));
MQQ1068:ROM32_INSTR_PT(107) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110100"));
MQQ1069:ROM32_INSTR_PT(108) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001001100"));
MQQ1070:ROM32_INSTR_PT(109) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001001100"));
MQQ1071:ROM32_INSTR_PT(110) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001100"));
MQQ1072:ROM32_INSTR_PT(111) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001100"));
MQQ1073:ROM32_INSTR_PT(112) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001100"));
MQQ1074:ROM32_INSTR_PT(113) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101100"));
MQQ1075:ROM32_INSTR_PT(114) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100101100"));
MQQ1076:ROM32_INSTR_PT(115) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010101100"));
MQQ1077:ROM32_INSTR_PT(116) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101100"));
MQQ1078:ROM32_INSTR_PT(117) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101100"));
MQQ1079:ROM32_INSTR_PT(118) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ1080:ROM32_INSTR_PT(119) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ1081:ROM32_INSTR_PT(120) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011100"));
MQQ1082:ROM32_INSTR_PT(121) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011100"));
MQQ1083:ROM32_INSTR_PT(122) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011011100"));
MQQ1084:ROM32_INSTR_PT(123) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ1085:ROM32_INSTR_PT(124) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111100"));
MQQ1086:ROM32_INSTR_PT(125) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ1087:ROM32_INSTR_PT(126) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ1088:ROM32_INSTR_PT(127) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011100"));
MQQ1089:ROM32_INSTR_PT(128) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111100"));
MQQ1090:ROM32_INSTR_PT(129) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ1091:ROM32_INSTR_PT(130) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ1092:ROM32_INSTR_PT(131) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001100"));
MQQ1093:ROM32_INSTR_PT(132) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101100"));
MQQ1094:ROM32_INSTR_PT(133) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ1095:ROM32_INSTR_PT(134) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111100"));
MQQ1096:ROM32_INSTR_PT(135) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111100"));
MQQ1097:ROM32_INSTR_PT(136) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011100"));
MQQ1098:ROM32_INSTR_PT(137) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0100100"));
MQQ1099:ROM32_INSTR_PT(138) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010100"));
MQQ1100:ROM32_INSTR_PT(139) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010100"));
MQQ1101:ROM32_INSTR_PT(140) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001100"));
MQQ1102:ROM32_INSTR_PT(141) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001100"));
MQQ1103:ROM32_INSTR_PT(142) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ1104:ROM32_INSTR_PT(143) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011100"));
MQQ1105:ROM32_INSTR_PT(144) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ1106:ROM32_INSTR_PT(145) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101100"));
MQQ1107:ROM32_INSTR_PT(146) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001100"));
MQQ1108:ROM32_INSTR_PT(147) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000000"));
MQQ1109:ROM32_INSTR_PT(148) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010000"));
MQQ1110:ROM32_INSTR_PT(149) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010000"));
MQQ1111:ROM32_INSTR_PT(150) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001000"));
MQQ1112:ROM32_INSTR_PT(151) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001000"));
MQQ1113:ROM32_INSTR_PT(152) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1000"));
MQQ1114:ROM32_INSTR_PT(153) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000100"));
MQQ1115:ROM32_INSTR_PT(154) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000100"));
MQQ1116:ROM32_INSTR_PT(155) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100100"));
MQQ1117:ROM32_INSTR_PT(156) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("00100"));
MQQ1118:ROM32_INSTR_PT(157) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010100"));
MQQ1119:ROM32_INSTR_PT(158) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111100"));
MQQ1120:ROM32_INSTR_PT(159) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111100"));
MQQ1121:ROM32_INSTR_PT(160) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011100"));
MQQ1122:ROM32_INSTR_PT(161) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111100"));
MQQ1123:ROM32_INSTR_PT(162) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011100"));
MQQ1124:ROM32_INSTR_PT(163) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111100"));
MQQ1125:ROM32_INSTR_PT(164) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000100"));
MQQ1126:ROM32_INSTR_PT(165) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101100"));
MQQ1127:ROM32_INSTR_PT(166) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ1128:ROM32_INSTR_PT(167) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("01100"));
MQQ1129:ROM32_INSTR_PT(168) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("10100"));
MQQ1130:ROM32_INSTR_PT(169) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000010"));
MQQ1131:ROM32_INSTR_PT(170) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000010"));
MQQ1132:ROM32_INSTR_PT(171) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000010"));
MQQ1133:ROM32_INSTR_PT(172) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000010"));
MQQ1134:ROM32_INSTR_PT(173) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100010"));
MQQ1135:ROM32_INSTR_PT(174) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100010"));
MQQ1136:ROM32_INSTR_PT(175) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000010"));
MQQ1137:ROM32_INSTR_PT(176) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ1138:ROM32_INSTR_PT(177) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010010"));
MQQ1139:ROM32_INSTR_PT(178) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110010"));
MQQ1140:ROM32_INSTR_PT(179) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001110010"));
MQQ1141:ROM32_INSTR_PT(180) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110010"));
MQQ1142:ROM32_INSTR_PT(181) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ1143:ROM32_INSTR_PT(182) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010010"));
MQQ1144:ROM32_INSTR_PT(183) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010010"));
MQQ1145:ROM32_INSTR_PT(184) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110010"));
MQQ1146:ROM32_INSTR_PT(185) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110010"));
MQQ1147:ROM32_INSTR_PT(186) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ1148:ROM32_INSTR_PT(187) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000010"));
MQQ1149:ROM32_INSTR_PT(188) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000010"));
MQQ1150:ROM32_INSTR_PT(189) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100010"));
MQQ1151:ROM32_INSTR_PT(190) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ1152:ROM32_INSTR_PT(191) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("000010"));
MQQ1153:ROM32_INSTR_PT(192) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010010"));
MQQ1154:ROM32_INSTR_PT(193) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110010"));
MQQ1155:ROM32_INSTR_PT(194) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110010"));
MQQ1156:ROM32_INSTR_PT(195) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110010"));
MQQ1157:ROM32_INSTR_PT(196) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ1158:ROM32_INSTR_PT(197) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110010"));
MQQ1159:ROM32_INSTR_PT(198) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ1160:ROM32_INSTR_PT(199) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001010"));
MQQ1161:ROM32_INSTR_PT(200) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001010"));
MQQ1162:ROM32_INSTR_PT(201) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101001010"));
MQQ1163:ROM32_INSTR_PT(202) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001001010"));
MQQ1164:ROM32_INSTR_PT(203) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001010"));
MQQ1165:ROM32_INSTR_PT(204) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001010"));
MQQ1166:ROM32_INSTR_PT(205) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100101010"));
MQQ1167:ROM32_INSTR_PT(206) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101010"));
MQQ1168:ROM32_INSTR_PT(207) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101010"));
MQQ1169:ROM32_INSTR_PT(208) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101010"));
MQQ1170:ROM32_INSTR_PT(209) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101010"));
MQQ1171:ROM32_INSTR_PT(210) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101010"));
MQQ1172:ROM32_INSTR_PT(211) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001010"));
MQQ1173:ROM32_INSTR_PT(212) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011010"));
MQQ1174:ROM32_INSTR_PT(213) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ1175:ROM32_INSTR_PT(214) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011010"));
MQQ1176:ROM32_INSTR_PT(215) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011011010"));
MQQ1177:ROM32_INSTR_PT(216) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111010"));
MQQ1178:ROM32_INSTR_PT(217) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111010"));
MQQ1179:ROM32_INSTR_PT(218) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011111010"));
MQQ1180:ROM32_INSTR_PT(219) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111010"));
MQQ1181:ROM32_INSTR_PT(220) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111010"));
MQQ1182:ROM32_INSTR_PT(221) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011010"));
MQQ1183:ROM32_INSTR_PT(222) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100111010"));
MQQ1184:ROM32_INSTR_PT(223) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111010"));
MQQ1185:ROM32_INSTR_PT(224) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111010"));
MQQ1186:ROM32_INSTR_PT(225) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101010"));
MQQ1187:ROM32_INSTR_PT(226) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011010"));
MQQ1188:ROM32_INSTR_PT(227) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ1189:ROM32_INSTR_PT(228) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100010"));
MQQ1190:ROM32_INSTR_PT(229) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100010"));
MQQ1191:ROM32_INSTR_PT(230) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ1192:ROM32_INSTR_PT(231) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001010"));
MQQ1193:ROM32_INSTR_PT(232) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001010"));
MQQ1194:ROM32_INSTR_PT(233) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101010"));
MQQ1195:ROM32_INSTR_PT(234) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011010"));
MQQ1196:ROM32_INSTR_PT(235) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011010"));
MQQ1197:ROM32_INSTR_PT(236) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011010"));
MQQ1198:ROM32_INSTR_PT(237) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110000110"));
MQQ1199:ROM32_INSTR_PT(238) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000110"));
MQQ1200:ROM32_INSTR_PT(239) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000110"));
MQQ1201:ROM32_INSTR_PT(240) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000110"));
MQQ1202:ROM32_INSTR_PT(241) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000110"));
MQQ1203:ROM32_INSTR_PT(242) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111000110"));
MQQ1204:ROM32_INSTR_PT(243) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000110"));
MQQ1205:ROM32_INSTR_PT(244) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000100110"));
MQQ1206:ROM32_INSTR_PT(245) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001100110"));
MQQ1207:ROM32_INSTR_PT(246) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000110"));
MQQ1208:ROM32_INSTR_PT(247) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000110"));
MQQ1209:ROM32_INSTR_PT(248) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100110"));
MQQ1210:ROM32_INSTR_PT(249) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100110"));
MQQ1211:ROM32_INSTR_PT(250) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110010110"));
MQQ1212:ROM32_INSTR_PT(251) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010110"));
MQQ1213:ROM32_INSTR_PT(252) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010110"));
MQQ1214:ROM32_INSTR_PT(253) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110110"));
MQQ1215:ROM32_INSTR_PT(254) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110110"));
MQQ1216:ROM32_INSTR_PT(255) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100110110"));
MQQ1217:ROM32_INSTR_PT(256) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110110"));
MQQ1218:ROM32_INSTR_PT(257) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110110"));
MQQ1219:ROM32_INSTR_PT(258) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100110"));
MQQ1220:ROM32_INSTR_PT(259) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010110"));
MQQ1221:ROM32_INSTR_PT(260) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100110110"));
MQQ1222:ROM32_INSTR_PT(261) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110110"));
MQQ1223:ROM32_INSTR_PT(262) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110110"));
MQQ1224:ROM32_INSTR_PT(263) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010110"));
MQQ1225:ROM32_INSTR_PT(264) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100001110"));
MQQ1226:ROM32_INSTR_PT(265) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001110"));
MQQ1227:ROM32_INSTR_PT(266) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110001110"));
MQQ1228:ROM32_INSTR_PT(267) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001110"));
MQQ1229:ROM32_INSTR_PT(268) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001110"));
MQQ1230:ROM32_INSTR_PT(269) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000101110"));
MQQ1231:ROM32_INSTR_PT(270) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100101110"));
MQQ1232:ROM32_INSTR_PT(271) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101110"));
MQQ1233:ROM32_INSTR_PT(272) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101110"));
MQQ1234:ROM32_INSTR_PT(273) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101110"));
MQQ1235:ROM32_INSTR_PT(274) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101110"));
MQQ1236:ROM32_INSTR_PT(275) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011110"));
MQQ1237:ROM32_INSTR_PT(276) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011110"));
MQQ1238:ROM32_INSTR_PT(277) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ1239:ROM32_INSTR_PT(278) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111110"));
MQQ1240:ROM32_INSTR_PT(279) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111110"));
MQQ1241:ROM32_INSTR_PT(280) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111110"));
MQQ1242:ROM32_INSTR_PT(281) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011110"));
MQQ1243:ROM32_INSTR_PT(282) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ1244:ROM32_INSTR_PT(283) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111110"));
MQQ1245:ROM32_INSTR_PT(284) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111110"));
MQQ1246:ROM32_INSTR_PT(285) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111110"));
MQQ1247:ROM32_INSTR_PT(286) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111110"));
MQQ1248:ROM32_INSTR_PT(287) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111110"));
MQQ1249:ROM32_INSTR_PT(288) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ1250:ROM32_INSTR_PT(289) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110110"));
MQQ1251:ROM32_INSTR_PT(290) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110110"));
MQQ1252:ROM32_INSTR_PT(291) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100110"));
MQQ1253:ROM32_INSTR_PT(292) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001110"));
MQQ1254:ROM32_INSTR_PT(293) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ1255:ROM32_INSTR_PT(294) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011110"));
MQQ1256:ROM32_INSTR_PT(295) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111110"));
MQQ1257:ROM32_INSTR_PT(296) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101110"));
MQQ1258:ROM32_INSTR_PT(297) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011110"));
MQQ1259:ROM32_INSTR_PT(298) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ1260:ROM32_INSTR_PT(299) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101110"));
MQQ1261:ROM32_INSTR_PT(300) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000010"));
MQQ1262:ROM32_INSTR_PT(301) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ1263:ROM32_INSTR_PT(302) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011010"));
MQQ1264:ROM32_INSTR_PT(303) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ1265:ROM32_INSTR_PT(304) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011010"));
MQQ1266:ROM32_INSTR_PT(305) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101010"));
MQQ1267:ROM32_INSTR_PT(306) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000110"));
MQQ1268:ROM32_INSTR_PT(307) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000110"));
MQQ1269:ROM32_INSTR_PT(308) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010110"));
MQQ1270:ROM32_INSTR_PT(309) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110110"));
MQQ1271:ROM32_INSTR_PT(310) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001110"));
MQQ1272:ROM32_INSTR_PT(311) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001110"));
MQQ1273:ROM32_INSTR_PT(312) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111110"));
MQQ1274:ROM32_INSTR_PT(313) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ1275:ROM32_INSTR_PT(314) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010110"));
MQQ1276:ROM32_INSTR_PT(315) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101110"));
MQQ1277:ROM32_INSTR_PT(316) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010010"));
MQQ1278:ROM32_INSTR_PT(317) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011010"));
MQQ1279:ROM32_INSTR_PT(318) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ1280:ROM32_INSTR_PT(319) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0000010"));
MQQ1281:ROM32_INSTR_PT(320) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000000"));
MQQ1282:ROM32_INSTR_PT(321) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010000"));
MQQ1283:ROM32_INSTR_PT(322) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101000"));
MQQ1284:ROM32_INSTR_PT(323) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101000"));
MQQ1285:ROM32_INSTR_PT(324) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101000"));
MQQ1286:ROM32_INSTR_PT(325) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100000"));
MQQ1287:ROM32_INSTR_PT(326) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0000100"));
MQQ1288:ROM32_INSTR_PT(327) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000100"));
MQQ1289:ROM32_INSTR_PT(328) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000100"));
MQQ1290:ROM32_INSTR_PT(329) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000100"));
MQQ1291:ROM32_INSTR_PT(330) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0100100"));
MQQ1292:ROM32_INSTR_PT(331) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001100"));
MQQ1293:ROM32_INSTR_PT(332) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00101100"));
MQQ1294:ROM32_INSTR_PT(333) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011100"));
MQQ1295:ROM32_INSTR_PT(334) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000000"));
MQQ1296:ROM32_INSTR_PT(335) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ1297:ROM32_INSTR_PT(336) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100010"));
MQQ1298:ROM32_INSTR_PT(337) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010010"));
MQQ1299:ROM32_INSTR_PT(338) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110010"));
MQQ1300:ROM32_INSTR_PT(339) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ1301:ROM32_INSTR_PT(340) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001010"));
MQQ1302:ROM32_INSTR_PT(341) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001010"));
MQQ1303:ROM32_INSTR_PT(342) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100110"));
MQQ1304:ROM32_INSTR_PT(343) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ1305:ROM32_INSTR_PT(344) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ1306:ROM32_INSTR_PT(345) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101110"));
MQQ1307:ROM32_INSTR_PT(346) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ1308:ROM32_INSTR_PT(347) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011110"));
MQQ1309:ROM32_INSTR_PT(348) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011110"));
MQQ1310:ROM32_INSTR_PT(349) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100110"));
MQQ1311:ROM32_INSTR_PT(350) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011110"));
MQQ1312:ROM32_INSTR_PT(351) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000000"));
MQQ1313:ROM32_INSTR_PT(352) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101000"));
MQQ1314:ROM32_INSTR_PT(353) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ1315:ROM32_INSTR_PT(354) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000010"));
MQQ1316:ROM32_INSTR_PT(355) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100010"));
MQQ1317:ROM32_INSTR_PT(356) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110110"));
MQQ1318:ROM32_INSTR_PT(357) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011110"));
MQQ1319:ROM32_INSTR_PT(358) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100010"));
MQQ1320:ROM32_INSTR_PT(359) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000001"));
MQQ1321:ROM32_INSTR_PT(360) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000001"));
MQQ1322:ROM32_INSTR_PT(361) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110000001"));
MQQ1323:ROM32_INSTR_PT(362) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000001"));
MQQ1324:ROM32_INSTR_PT(363) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100001"));
MQQ1325:ROM32_INSTR_PT(364) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11100001"));
MQQ1326:ROM32_INSTR_PT(365) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000001"));
MQQ1327:ROM32_INSTR_PT(366) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ1328:ROM32_INSTR_PT(367) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010001"));
MQQ1329:ROM32_INSTR_PT(368) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010001"));
MQQ1330:ROM32_INSTR_PT(369) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110001"));
MQQ1331:ROM32_INSTR_PT(370) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110001"));
MQQ1332:ROM32_INSTR_PT(371) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001110001"));
MQQ1333:ROM32_INSTR_PT(372) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00110001"));
MQQ1334:ROM32_INSTR_PT(373) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110001"));
MQQ1335:ROM32_INSTR_PT(374) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110001"));
MQQ1336:ROM32_INSTR_PT(375) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110001"));
MQQ1337:ROM32_INSTR_PT(376) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110001"));
MQQ1338:ROM32_INSTR_PT(377) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110001"));
MQQ1339:ROM32_INSTR_PT(378) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000001"));
MQQ1340:ROM32_INSTR_PT(379) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ1341:ROM32_INSTR_PT(380) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0100001"));
MQQ1342:ROM32_INSTR_PT(381) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100001"));
MQQ1343:ROM32_INSTR_PT(382) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010001"));
MQQ1344:ROM32_INSTR_PT(383) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100110001"));
MQQ1345:ROM32_INSTR_PT(384) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110001"));
MQQ1346:ROM32_INSTR_PT(385) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010001"));
MQQ1347:ROM32_INSTR_PT(386) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001001"));
MQQ1348:ROM32_INSTR_PT(387) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001001"));
MQQ1349:ROM32_INSTR_PT(388) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111001001"));
MQQ1350:ROM32_INSTR_PT(389) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001001"));
MQQ1351:ROM32_INSTR_PT(390) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001001"));
MQQ1352:ROM32_INSTR_PT(391) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101001"));
MQQ1353:ROM32_INSTR_PT(392) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100101001"));
MQQ1354:ROM32_INSTR_PT(393) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101001"));
MQQ1355:ROM32_INSTR_PT(394) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001101001"));
MQQ1356:ROM32_INSTR_PT(395) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101001"));
MQQ1357:ROM32_INSTR_PT(396) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101001"));
MQQ1358:ROM32_INSTR_PT(397) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111101001"));
MQQ1359:ROM32_INSTR_PT(398) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110011001"));
MQQ1360:ROM32_INSTR_PT(399) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001011001"));
MQQ1361:ROM32_INSTR_PT(400) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011111001"));
MQQ1362:ROM32_INSTR_PT(401) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111001"));
MQQ1363:ROM32_INSTR_PT(402) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011001"));
MQQ1364:ROM32_INSTR_PT(403) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011001"));
MQQ1365:ROM32_INSTR_PT(404) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111001"));
MQQ1366:ROM32_INSTR_PT(405) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111001"));
MQQ1367:ROM32_INSTR_PT(406) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111001"));
MQQ1368:ROM32_INSTR_PT(407) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011001"));
MQQ1369:ROM32_INSTR_PT(408) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110111001"));
MQQ1370:ROM32_INSTR_PT(409) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111001"));
MQQ1371:ROM32_INSTR_PT(410) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011001"));
MQQ1372:ROM32_INSTR_PT(411) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000001"));
MQQ1373:ROM32_INSTR_PT(412) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ1374:ROM32_INSTR_PT(413) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100001"));
MQQ1375:ROM32_INSTR_PT(414) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0010001"));
MQQ1376:ROM32_INSTR_PT(415) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010001"));
MQQ1377:ROM32_INSTR_PT(416) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001001"));
MQQ1378:ROM32_INSTR_PT(417) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101001"));
MQQ1379:ROM32_INSTR_PT(418) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011001"));
MQQ1380:ROM32_INSTR_PT(419) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011001"));
MQQ1381:ROM32_INSTR_PT(420) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000101"));
MQQ1382:ROM32_INSTR_PT(421) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101000101"));
MQQ1383:ROM32_INSTR_PT(422) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000101"));
MQQ1384:ROM32_INSTR_PT(423) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000101"));
MQQ1385:ROM32_INSTR_PT(424) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000101"));
MQQ1386:ROM32_INSTR_PT(425) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000101"));
MQQ1387:ROM32_INSTR_PT(426) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100101"));
MQQ1388:ROM32_INSTR_PT(427) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100101"));
MQQ1389:ROM32_INSTR_PT(428) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001100101"));
MQQ1390:ROM32_INSTR_PT(429) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001100101"));
MQQ1391:ROM32_INSTR_PT(430) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100101"));
MQQ1392:ROM32_INSTR_PT(431) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11100101"));
MQQ1393:ROM32_INSTR_PT(432) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100101"));
MQQ1394:ROM32_INSTR_PT(433) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110010101"));
MQQ1395:ROM32_INSTR_PT(434) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001010101"));
MQQ1396:ROM32_INSTR_PT(435) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101010101"));
MQQ1397:ROM32_INSTR_PT(436) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010101"));
MQQ1398:ROM32_INSTR_PT(437) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110101"));
MQQ1399:ROM32_INSTR_PT(438) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110101"));
MQQ1400:ROM32_INSTR_PT(439) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110101"));
MQQ1401:ROM32_INSTR_PT(440) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110101"));
MQQ1402:ROM32_INSTR_PT(441) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110101"));
MQQ1403:ROM32_INSTR_PT(442) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000101"));
MQQ1404:ROM32_INSTR_PT(443) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000101"));
MQQ1405:ROM32_INSTR_PT(444) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100101"));
MQQ1406:ROM32_INSTR_PT(445) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010101"));
MQQ1407:ROM32_INSTR_PT(446) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110101"));
MQQ1408:ROM32_INSTR_PT(447) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110101"));
MQQ1409:ROM32_INSTR_PT(448) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010101"));
MQQ1410:ROM32_INSTR_PT(449) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0100001101"));
MQQ1411:ROM32_INSTR_PT(450) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110001101"));
MQQ1412:ROM32_INSTR_PT(451) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001001101"));
MQQ1413:ROM32_INSTR_PT(452) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011001101"));
MQQ1414:ROM32_INSTR_PT(453) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101101"));
MQQ1415:ROM32_INSTR_PT(454) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101101"));
MQQ1416:ROM32_INSTR_PT(455) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001101"));
MQQ1417:ROM32_INSTR_PT(456) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001101"));
MQQ1418:ROM32_INSTR_PT(457) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101101"));
MQQ1419:ROM32_INSTR_PT(458) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101101"));
MQQ1420:ROM32_INSTR_PT(459) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011101"));
MQQ1421:ROM32_INSTR_PT(460) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011101"));
MQQ1422:ROM32_INSTR_PT(461) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111101"));
MQQ1423:ROM32_INSTR_PT(462) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011101"));
MQQ1424:ROM32_INSTR_PT(463) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011101"));
MQQ1425:ROM32_INSTR_PT(464) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111101"));
MQQ1426:ROM32_INSTR_PT(465) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("100111101"));
MQQ1427:ROM32_INSTR_PT(466) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111101"));
MQQ1428:ROM32_INSTR_PT(467) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111101"));
MQQ1429:ROM32_INSTR_PT(468) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100101"));
MQQ1430:ROM32_INSTR_PT(469) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010101"));
MQQ1431:ROM32_INSTR_PT(470) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0010101"));
MQQ1432:ROM32_INSTR_PT(471) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110101"));
MQQ1433:ROM32_INSTR_PT(472) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010101"));
MQQ1434:ROM32_INSTR_PT(473) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001101"));
MQQ1435:ROM32_INSTR_PT(474) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001101"));
MQQ1436:ROM32_INSTR_PT(475) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001101"));
MQQ1437:ROM32_INSTR_PT(476) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011101"));
MQQ1438:ROM32_INSTR_PT(477) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011101"));
MQQ1439:ROM32_INSTR_PT(478) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111101"));
MQQ1440:ROM32_INSTR_PT(479) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ1441:ROM32_INSTR_PT(480) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010001"));
MQQ1442:ROM32_INSTR_PT(481) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110001"));
MQQ1443:ROM32_INSTR_PT(482) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001001"));
MQQ1444:ROM32_INSTR_PT(483) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101001"));
MQQ1445:ROM32_INSTR_PT(484) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011001"));
MQQ1446:ROM32_INSTR_PT(485) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111001"));
MQQ1447:ROM32_INSTR_PT(486) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111001"));
MQQ1448:ROM32_INSTR_PT(487) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011001"));
MQQ1449:ROM32_INSTR_PT(488) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011001"));
MQQ1450:ROM32_INSTR_PT(489) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000101"));
MQQ1451:ROM32_INSTR_PT(490) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100101"));
MQQ1452:ROM32_INSTR_PT(491) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11010101"));
MQQ1453:ROM32_INSTR_PT(492) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100101"));
MQQ1454:ROM32_INSTR_PT(493) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010101"));
MQQ1455:ROM32_INSTR_PT(494) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111101"));
MQQ1456:ROM32_INSTR_PT(495) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011101"));
MQQ1457:ROM32_INSTR_PT(496) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111101"));
MQQ1458:ROM32_INSTR_PT(497) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101101"));
MQQ1459:ROM32_INSTR_PT(498) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001101"));
MQQ1460:ROM32_INSTR_PT(499) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0000001"));
MQQ1461:ROM32_INSTR_PT(500) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001"));
MQQ1462:ROM32_INSTR_PT(501) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000011"));
MQQ1463:ROM32_INSTR_PT(502) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101000011"));
MQQ1464:ROM32_INSTR_PT(503) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000011"));
MQQ1465:ROM32_INSTR_PT(504) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000011"));
MQQ1466:ROM32_INSTR_PT(505) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010100011"));
MQQ1467:ROM32_INSTR_PT(506) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100011"));
MQQ1468:ROM32_INSTR_PT(507) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100011"));
MQQ1469:ROM32_INSTR_PT(508) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000000011"));
MQQ1470:ROM32_INSTR_PT(509) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100011"));
MQQ1471:ROM32_INSTR_PT(510) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000011"));
MQQ1472:ROM32_INSTR_PT(511) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010011"));
MQQ1473:ROM32_INSTR_PT(512) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010010011"));
MQQ1474:ROM32_INSTR_PT(513) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010011"));
MQQ1475:ROM32_INSTR_PT(514) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010011"));
MQQ1476:ROM32_INSTR_PT(515) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010011"));
MQQ1477:ROM32_INSTR_PT(516) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("101110011"));
MQQ1478:ROM32_INSTR_PT(517) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001110011"));
MQQ1479:ROM32_INSTR_PT(518) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00010011"));
MQQ1480:ROM32_INSTR_PT(519) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110011"));
MQQ1481:ROM32_INSTR_PT(520) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110011"));
MQQ1482:ROM32_INSTR_PT(521) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110011"));
MQQ1483:ROM32_INSTR_PT(522) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000011"));
MQQ1484:ROM32_INSTR_PT(523) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000011"));
MQQ1485:ROM32_INSTR_PT(524) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100011"));
MQQ1486:ROM32_INSTR_PT(525) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ1487:ROM32_INSTR_PT(526) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1100011"));
MQQ1488:ROM32_INSTR_PT(527) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010011"));
MQQ1489:ROM32_INSTR_PT(528) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000110011"));
MQQ1490:ROM32_INSTR_PT(529) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1010011"));
MQQ1491:ROM32_INSTR_PT(530) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001011"));
MQQ1492:ROM32_INSTR_PT(531) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101001011"));
MQQ1493:ROM32_INSTR_PT(532) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001001011"));
MQQ1494:ROM32_INSTR_PT(533) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("111001011"));
MQQ1495:ROM32_INSTR_PT(534) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0000101011"));
MQQ1496:ROM32_INSTR_PT(535) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110101011"));
MQQ1497:ROM32_INSTR_PT(536) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011101011"));
MQQ1498:ROM32_INSTR_PT(537) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101011"));
MQQ1499:ROM32_INSTR_PT(538) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101011"));
MQQ1500:ROM32_INSTR_PT(539) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101011"));
MQQ1501:ROM32_INSTR_PT(540) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011011"));
MQQ1502:ROM32_INSTR_PT(541) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ1503:ROM32_INSTR_PT(542) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011011"));
MQQ1504:ROM32_INSTR_PT(543) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111011"));
MQQ1505:ROM32_INSTR_PT(544) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011011"));
MQQ1506:ROM32_INSTR_PT(545) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ1507:ROM32_INSTR_PT(546) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111011"));
MQQ1508:ROM32_INSTR_PT(547) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101011"));
MQQ1509:ROM32_INSTR_PT(548) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011011"));
MQQ1510:ROM32_INSTR_PT(549) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111011"));
MQQ1511:ROM32_INSTR_PT(550) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100011"));
MQQ1512:ROM32_INSTR_PT(551) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100011"));
MQQ1513:ROM32_INSTR_PT(552) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10110011"));
MQQ1514:ROM32_INSTR_PT(553) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00001011"));
MQQ1515:ROM32_INSTR_PT(554) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001011"));
MQQ1516:ROM32_INSTR_PT(555) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1101011"));
MQQ1517:ROM32_INSTR_PT(556) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000011011"));
MQQ1518:ROM32_INSTR_PT(557) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011011"));
MQQ1519:ROM32_INSTR_PT(558) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011011"));
MQQ1520:ROM32_INSTR_PT(559) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111011"));
MQQ1521:ROM32_INSTR_PT(560) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101011"));
MQQ1522:ROM32_INSTR_PT(561) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0011011"));
MQQ1523:ROM32_INSTR_PT(562) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111011"));
MQQ1524:ROM32_INSTR_PT(563) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111011"));
MQQ1525:ROM32_INSTR_PT(564) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ1526:ROM32_INSTR_PT(565) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000111"));
MQQ1527:ROM32_INSTR_PT(566) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000111"));
MQQ1528:ROM32_INSTR_PT(567) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000111"));
MQQ1529:ROM32_INSTR_PT(568) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001000111"));
MQQ1530:ROM32_INSTR_PT(569) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000111"));
MQQ1531:ROM32_INSTR_PT(570) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011000111"));
MQQ1532:ROM32_INSTR_PT(571) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010100111"));
MQQ1533:ROM32_INSTR_PT(572) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100111"));
MQQ1534:ROM32_INSTR_PT(573) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10100111"));
MQQ1535:ROM32_INSTR_PT(574) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001100111"));
MQQ1536:ROM32_INSTR_PT(575) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011100111"));
MQQ1537:ROM32_INSTR_PT(576) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000111"));
MQQ1538:ROM32_INSTR_PT(577) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000111"));
MQQ1539:ROM32_INSTR_PT(578) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000010111"));
MQQ1540:ROM32_INSTR_PT(579) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010111"));
MQQ1541:ROM32_INSTR_PT(580) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001010111"));
MQQ1542:ROM32_INSTR_PT(581) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("011010111"));
MQQ1543:ROM32_INSTR_PT(582) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110110111"));
MQQ1544:ROM32_INSTR_PT(583) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010111"));
MQQ1545:ROM32_INSTR_PT(584) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01100111"));
MQQ1546:ROM32_INSTR_PT(585) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000001111"));
MQQ1547:ROM32_INSTR_PT(586) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010001111"));
MQQ1548:ROM32_INSTR_PT(587) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001111"));
MQQ1549:ROM32_INSTR_PT(588) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001111"));
MQQ1550:ROM32_INSTR_PT(589) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001111"));
MQQ1551:ROM32_INSTR_PT(590) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000101111"));
MQQ1552:ROM32_INSTR_PT(591) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0001101111"));
MQQ1553:ROM32_INSTR_PT(592) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101111"));
MQQ1554:ROM32_INSTR_PT(593) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101111"));
MQQ1555:ROM32_INSTR_PT(594) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0001111"));
MQQ1556:ROM32_INSTR_PT(595) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11101111"));
MQQ1557:ROM32_INSTR_PT(596) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011111"));
MQQ1558:ROM32_INSTR_PT(597) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011111"));
MQQ1559:ROM32_INSTR_PT(598) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("001011111"));
MQQ1560:ROM32_INSTR_PT(599) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111111"));
MQQ1561:ROM32_INSTR_PT(600) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111111"));
MQQ1562:ROM32_INSTR_PT(601) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ1563:ROM32_INSTR_PT(602) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011111"));
MQQ1564:ROM32_INSTR_PT(603) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ1565:ROM32_INSTR_PT(604) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111111"));
MQQ1566:ROM32_INSTR_PT(605) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111111"));
MQQ1567:ROM32_INSTR_PT(606) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11111111"));
MQQ1568:ROM32_INSTR_PT(607) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01101111"));
MQQ1569:ROM32_INSTR_PT(608) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ1570:ROM32_INSTR_PT(609) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10111111"));
MQQ1571:ROM32_INSTR_PT(610) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111111"));
MQQ1572:ROM32_INSTR_PT(611) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1573:ROM32_INSTR_PT(612) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1574:ROM32_INSTR_PT(613) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000111"));
MQQ1575:ROM32_INSTR_PT(614) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110111"));
MQQ1576:ROM32_INSTR_PT(615) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110111"));
MQQ1577:ROM32_INSTR_PT(616) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000111"));
MQQ1578:ROM32_INSTR_PT(617) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001111"));
MQQ1579:ROM32_INSTR_PT(618) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011111"));
MQQ1580:ROM32_INSTR_PT(619) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ1581:ROM32_INSTR_PT(620) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01011111"));
MQQ1582:ROM32_INSTR_PT(621) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01111111"));
MQQ1583:ROM32_INSTR_PT(622) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ1584:ROM32_INSTR_PT(623) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ1585:ROM32_INSTR_PT(624) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ1586:ROM32_INSTR_PT(625) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ1587:ROM32_INSTR_PT(626) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ1588:ROM32_INSTR_PT(627) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000011"));
MQQ1589:ROM32_INSTR_PT(628) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("10011"));
MQQ1590:ROM32_INSTR_PT(629) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ1591:ROM32_INSTR_PT(630) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011011"));
MQQ1592:ROM32_INSTR_PT(631) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000111011"));
MQQ1593:ROM32_INSTR_PT(632) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00111011"));
MQQ1594:ROM32_INSTR_PT(633) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111011"));
MQQ1595:ROM32_INSTR_PT(634) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ1596:ROM32_INSTR_PT(635) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ1597:ROM32_INSTR_PT(636) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011011"));
MQQ1598:ROM32_INSTR_PT(637) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("10011"));
MQQ1599:ROM32_INSTR_PT(638) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("010000111"));
MQQ1600:ROM32_INSTR_PT(639) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100111"));
MQQ1601:ROM32_INSTR_PT(640) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010111"));
MQQ1602:ROM32_INSTR_PT(641) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000111"));
MQQ1603:ROM32_INSTR_PT(642) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ1604:ROM32_INSTR_PT(643) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1605:ROM32_INSTR_PT(644) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1606:ROM32_INSTR_PT(645) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0010111"));
MQQ1607:ROM32_INSTR_PT(646) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110111"));
MQQ1608:ROM32_INSTR_PT(647) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011111"));
MQQ1609:ROM32_INSTR_PT(648) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ1610:ROM32_INSTR_PT(649) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ1611:ROM32_INSTR_PT(650) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ1612:ROM32_INSTR_PT(651) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(8) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ1613:ROM32_INSTR_PT(652) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11000001"));
MQQ1614:ROM32_INSTR_PT(653) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000001"));
MQQ1615:ROM32_INSTR_PT(654) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110001"));
MQQ1616:ROM32_INSTR_PT(655) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110001"));
MQQ1617:ROM32_INSTR_PT(656) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001001"));
MQQ1618:ROM32_INSTR_PT(657) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101001"));
MQQ1619:ROM32_INSTR_PT(658) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001001"));
MQQ1620:ROM32_INSTR_PT(659) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00011001"));
MQQ1621:ROM32_INSTR_PT(660) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101001"));
MQQ1622:ROM32_INSTR_PT(661) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("00000101"));
MQQ1623:ROM32_INSTR_PT(662) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01000101"));
MQQ1624:ROM32_INSTR_PT(663) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("000100101"));
MQQ1625:ROM32_INSTR_PT(664) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11110101"));
MQQ1626:ROM32_INSTR_PT(665) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11001101"));
MQQ1627:ROM32_INSTR_PT(666) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011101"));
MQQ1628:ROM32_INSTR_PT(667) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011101"));
MQQ1629:ROM32_INSTR_PT(668) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000001"));
MQQ1630:ROM32_INSTR_PT(669) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011101"));
MQQ1631:ROM32_INSTR_PT(670) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("01001"));
MQQ1632:ROM32_INSTR_PT(671) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100101"));
MQQ1633:ROM32_INSTR_PT(672) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100011"));
MQQ1634:ROM32_INSTR_PT(673) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ1635:ROM32_INSTR_PT(674) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01110011"));
MQQ1636:ROM32_INSTR_PT(675) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("000011"));
MQQ1637:ROM32_INSTR_PT(676) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ1638:ROM32_INSTR_PT(677) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10101011"));
MQQ1639:ROM32_INSTR_PT(678) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10011011"));
MQQ1640:ROM32_INSTR_PT(679) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011011"));
MQQ1641:ROM32_INSTR_PT(680) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011011"));
MQQ1642:ROM32_INSTR_PT(681) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("010011"));
MQQ1643:ROM32_INSTR_PT(682) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("110100111"));
MQQ1644:ROM32_INSTR_PT(683) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10010111"));
MQQ1645:ROM32_INSTR_PT(684) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("01010111"));
MQQ1646:ROM32_INSTR_PT(685) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("10001111"));
MQQ1647:ROM32_INSTR_PT(686) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("101111"));
MQQ1648:ROM32_INSTR_PT(687) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011111"));
MQQ1649:ROM32_INSTR_PT(688) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ1650:ROM32_INSTR_PT(689) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0111111"));
MQQ1651:ROM32_INSTR_PT(690) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1652:ROM32_INSTR_PT(691) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000111"));
MQQ1653:ROM32_INSTR_PT(692) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1110111"));
MQQ1654:ROM32_INSTR_PT(693) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("11011111"));
MQQ1655:ROM32_INSTR_PT(694) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ1656:ROM32_INSTR_PT(695) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0011"));
MQQ1657:ROM32_INSTR_PT(696) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ1658:ROM32_INSTR_PT(697) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1659:ROM32_INSTR_PT(698) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0101111"));
MQQ1660:ROM32_INSTR_PT(699) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1011111"));
MQQ1661:ROM32_INSTR_PT(700) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ1662:ROM32_INSTR_PT(701) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("01111"));
MQQ1663:ROM32_INSTR_PT(702) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1000001"));
MQQ1664:ROM32_INSTR_PT(703) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1001001"));
MQQ1665:ROM32_INSTR_PT(704) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111001"));
MQQ1666:ROM32_INSTR_PT(705) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100001"));
MQQ1667:ROM32_INSTR_PT(706) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("001001"));
MQQ1668:ROM32_INSTR_PT(707) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111101"));
MQQ1669:ROM32_INSTR_PT(708) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("0110111"));
MQQ1670:ROM32_INSTR_PT(709) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1671:ROM32_INSTR_PT(710) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ1672:ROM32_INSTR_PT(711) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1673:ROM32_INSTR_PT(712) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100111"));
MQQ1674:ROM32_INSTR_PT(713) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("011111"));
MQQ1675:ROM32_INSTR_PT(714) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(9) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ1676:ROM32_INSTR_PT(715) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100101"));
MQQ1677:ROM32_INSTR_PT(716) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ1678:ROM32_INSTR_PT(717) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("0111"));
MQQ1679:ROM32_INSTR_PT(718) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(9)
     ) , STD_ULOGIC_VECTOR'("1101"));
MQQ1680:ROM32_INSTR_PT(719) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100000"));
MQQ1681:ROM32_INSTR_PT(720) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100000"));
MQQ1682:ROM32_INSTR_PT(721) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1010000"));
MQQ1683:ROM32_INSTR_PT(722) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000110000"));
MQQ1684:ROM32_INSTR_PT(723) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01110000"));
MQQ1685:ROM32_INSTR_PT(724) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100000"));
MQQ1686:ROM32_INSTR_PT(725) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111000"));
MQQ1687:ROM32_INSTR_PT(726) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0111000"));
MQQ1688:ROM32_INSTR_PT(727) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000100"));
MQQ1689:ROM32_INSTR_PT(728) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100100"));
MQQ1690:ROM32_INSTR_PT(729) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1100100"));
MQQ1691:ROM32_INSTR_PT(730) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1100100"));
MQQ1692:ROM32_INSTR_PT(731) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ1693:ROM32_INSTR_PT(732) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01101100"));
MQQ1694:ROM32_INSTR_PT(733) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("10011100"));
MQQ1695:ROM32_INSTR_PT(734) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101100"));
MQQ1696:ROM32_INSTR_PT(735) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01100"));
MQQ1697:ROM32_INSTR_PT(736) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100100"));
MQQ1698:ROM32_INSTR_PT(737) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100000"));
MQQ1699:ROM32_INSTR_PT(738) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1100000"));
MQQ1700:ROM32_INSTR_PT(739) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00000100"));
MQQ1701:ROM32_INSTR_PT(740) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0101100"));
MQQ1702:ROM32_INSTR_PT(741) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011100"));
MQQ1703:ROM32_INSTR_PT(742) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ1704:ROM32_INSTR_PT(743) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11100"));
MQQ1705:ROM32_INSTR_PT(744) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000"));
MQQ1706:ROM32_INSTR_PT(745) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01100010"));
MQQ1707:ROM32_INSTR_PT(746) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000010"));
MQQ1708:ROM32_INSTR_PT(747) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00010010"));
MQQ1709:ROM32_INSTR_PT(748) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00000010"));
MQQ1710:ROM32_INSTR_PT(749) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11001010"));
MQQ1711:ROM32_INSTR_PT(750) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111010"));
MQQ1712:ROM32_INSTR_PT(751) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01001010"));
MQQ1713:ROM32_INSTR_PT(752) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101010"));
MQQ1714:ROM32_INSTR_PT(753) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("010000110"));
MQQ1715:ROM32_INSTR_PT(754) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1000110"));
MQQ1716:ROM32_INSTR_PT(755) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("110100110"));
MQQ1717:ROM32_INSTR_PT(756) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0001110"));
MQQ1718:ROM32_INSTR_PT(757) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1001110"));
MQQ1719:ROM32_INSTR_PT(758) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011110"));
MQQ1720:ROM32_INSTR_PT(759) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("10011110"));
MQQ1721:ROM32_INSTR_PT(760) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1010010"));
MQQ1722:ROM32_INSTR_PT(761) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("0110"));
MQQ1723:ROM32_INSTR_PT(762) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011110"));
MQQ1724:ROM32_INSTR_PT(763) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1111110"));
MQQ1725:ROM32_INSTR_PT(764) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("010110"));
MQQ1726:ROM32_INSTR_PT(765) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("010100"));
MQQ1727:ROM32_INSTR_PT(766) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1101100"));
MQQ1728:ROM32_INSTR_PT(767) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011100"));
MQQ1729:ROM32_INSTR_PT(768) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110000"));
MQQ1730:ROM32_INSTR_PT(769) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("00100"));
MQQ1731:ROM32_INSTR_PT(770) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100010"));
MQQ1732:ROM32_INSTR_PT(771) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1001110"));
MQQ1733:ROM32_INSTR_PT(772) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("0000"));
MQQ1734:ROM32_INSTR_PT(773) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01110"));
MQQ1735:ROM32_INSTR_PT(774) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01000001"));
MQQ1736:ROM32_INSTR_PT(775) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("110100001"));
MQQ1737:ROM32_INSTR_PT(776) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01010001"));
MQQ1738:ROM32_INSTR_PT(777) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11010001"));
MQQ1739:ROM32_INSTR_PT(778) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1010001"));
MQQ1740:ROM32_INSTR_PT(779) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000001"));
MQQ1741:ROM32_INSTR_PT(780) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1000001"));
MQQ1742:ROM32_INSTR_PT(781) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("010001"));
MQQ1743:ROM32_INSTR_PT(782) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0001001"));
MQQ1744:ROM32_INSTR_PT(783) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("001001"));
MQQ1745:ROM32_INSTR_PT(784) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011001"));
MQQ1746:ROM32_INSTR_PT(785) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111001"));
MQQ1747:ROM32_INSTR_PT(786) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011001"));
MQQ1748:ROM32_INSTR_PT(787) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00100101"));
MQQ1749:ROM32_INSTR_PT(788) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00010101"));
MQQ1750:ROM32_INSTR_PT(789) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00011101"));
MQQ1751:ROM32_INSTR_PT(790) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("10011101"));
MQQ1752:ROM32_INSTR_PT(791) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011101"));
MQQ1753:ROM32_INSTR_PT(792) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110101"));
MQQ1754:ROM32_INSTR_PT(793) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("10101"));
MQQ1755:ROM32_INSTR_PT(794) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11101"));
MQQ1756:ROM32_INSTR_PT(795) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000101"));
MQQ1757:ROM32_INSTR_PT(796) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000101"));
MQQ1758:ROM32_INSTR_PT(797) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11101"));
MQQ1759:ROM32_INSTR_PT(798) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101101"));
MQQ1760:ROM32_INSTR_PT(799) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100001"));
MQQ1761:ROM32_INSTR_PT(800) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000100011"));
MQQ1762:ROM32_INSTR_PT(801) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00000011"));
MQQ1763:ROM32_INSTR_PT(802) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000011"));
MQQ1764:ROM32_INSTR_PT(803) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1010011"));
MQQ1765:ROM32_INSTR_PT(804) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("10011"));
MQQ1766:ROM32_INSTR_PT(805) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01001011"));
MQQ1767:ROM32_INSTR_PT(806) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0001011"));
MQQ1768:ROM32_INSTR_PT(807) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01000011"));
MQQ1769:ROM32_INSTR_PT(808) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101011"));
MQQ1770:ROM32_INSTR_PT(809) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ1771:ROM32_INSTR_PT(810) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100111"));
MQQ1772:ROM32_INSTR_PT(811) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("00010111"));
MQQ1773:ROM32_INSTR_PT(812) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01010111"));
MQQ1774:ROM32_INSTR_PT(813) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1775:ROM32_INSTR_PT(814) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1110111"));
MQQ1776:ROM32_INSTR_PT(815) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("11010111"));
MQQ1777:ROM32_INSTR_PT(816) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("000101111"));
MQQ1778:ROM32_INSTR_PT(817) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01101111"));
MQQ1779:ROM32_INSTR_PT(818) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1780:ROM32_INSTR_PT(819) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1781:ROM32_INSTR_PT(820) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ1782:ROM32_INSTR_PT(821) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1783:ROM32_INSTR_PT(822) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101011"));
MQQ1784:ROM32_INSTR_PT(823) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("01000111"));
MQQ1785:ROM32_INSTR_PT(824) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0110111"));
MQQ1786:ROM32_INSTR_PT(825) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1787:ROM32_INSTR_PT(826) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101111"));
MQQ1788:ROM32_INSTR_PT(827) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ1789:ROM32_INSTR_PT(828) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("0111"));
MQQ1790:ROM32_INSTR_PT(829) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1791:ROM32_INSTR_PT(830) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(7) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01111"));
MQQ1792:ROM32_INSTR_PT(831) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110001"));
MQQ1793:ROM32_INSTR_PT(832) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011001"));
MQQ1794:ROM32_INSTR_PT(833) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1001101"));
MQQ1795:ROM32_INSTR_PT(834) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("01001"));
MQQ1796:ROM32_INSTR_PT(835) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0100011"));
MQQ1797:ROM32_INSTR_PT(836) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1111011"));
MQQ1798:ROM32_INSTR_PT(837) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("11011"));
MQQ1799:ROM32_INSTR_PT(838) <=
    Eq(( ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("011"));
MQQ1800:ROM32_INSTR_PT(839) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("0000111"));
MQQ1801:ROM32_INSTR_PT(840) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("1111111"));
MQQ1802:ROM32_INSTR_PT(841) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011111"));
MQQ1803:ROM32_INSTR_PT(842) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("101111"));
MQQ1804:ROM32_INSTR_PT(843) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ1805:ROM32_INSTR_PT(844) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1806:ROM32_INSTR_PT(845) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("011111"));
MQQ1807:ROM32_INSTR_PT(846) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("000101"));
MQQ1808:ROM32_INSTR_PT(847) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("100011"));
MQQ1809:ROM32_INSTR_PT(848) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("1111"));
MQQ1810:ROM32_INSTR_PT(849) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(8) ) , STD_ULOGIC_VECTOR'("10111"));
MQQ1811:ROM32_INSTR_PT(850) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(8)
     ) , STD_ULOGIC_VECTOR'("0111"));
MQQ1812:ROM32_INSTR_PT(851) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1001000"));
MQQ1813:ROM32_INSTR_PT(852) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("110000"));
MQQ1814:ROM32_INSTR_PT(853) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("00011100"));
MQQ1815:ROM32_INSTR_PT(854) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("00000010"));
MQQ1816:ROM32_INSTR_PT(855) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0100010"));
MQQ1817:ROM32_INSTR_PT(856) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0000010"));
MQQ1818:ROM32_INSTR_PT(857) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("101110"));
MQQ1819:ROM32_INSTR_PT(858) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1101110"));
MQQ1820:ROM32_INSTR_PT(859) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1001100"));
MQQ1821:ROM32_INSTR_PT(860) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("00000"));
MQQ1822:ROM32_INSTR_PT(861) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("1110"));
MQQ1823:ROM32_INSTR_PT(862) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0100101"));
MQQ1824:ROM32_INSTR_PT(863) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1001101"));
MQQ1825:ROM32_INSTR_PT(864) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("001101"));
MQQ1826:ROM32_INSTR_PT(865) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1101101"));
MQQ1827:ROM32_INSTR_PT(866) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("1101"));
MQQ1828:ROM32_INSTR_PT(867) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1010011"));
MQQ1829:ROM32_INSTR_PT(868) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("1001011"));
MQQ1830:ROM32_INSTR_PT(869) <=
    Eq(( ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1831:ROM32_INSTR_PT(870) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("0011111"));
MQQ1832:ROM32_INSTR_PT(871) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("111111"));
MQQ1833:ROM32_INSTR_PT(872) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(6) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1834:ROM32_INSTR_PT(873) <=
    Eq(( ROM_ADDR_L2(1) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("11111"));
MQQ1835:ROM32_INSTR_PT(874) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6) & 
    ROM_ADDR_L2(7) ) , STD_ULOGIC_VECTOR'("01111"));
MQQ1836:ROM32_INSTR_PT(875) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("1101"));
MQQ1837:ROM32_INSTR_PT(876) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(7)
     ) , STD_ULOGIC_VECTOR'("000011"));
MQQ1838:ROM32_INSTR_PT(877) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) ) , STD_ULOGIC_VECTOR'("0000100"));
MQQ1839:ROM32_INSTR_PT(878) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(5) & ROM_ADDR_L2(6)
     ) , STD_ULOGIC_VECTOR'("010010"));
MQQ1840:ROM32_INSTR_PT(879) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(6)
     ) , STD_ULOGIC_VECTOR'("00"));
MQQ1841:ROM32_INSTR_PT(880) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5) & 
    ROM_ADDR_L2(6) ) , STD_ULOGIC_VECTOR'("111"));
MQQ1842:ROM32_INSTR_PT(881) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) & ROM_ADDR_L2(6)
     ) , STD_ULOGIC_VECTOR'("110111"));
MQQ1843:ROM32_INSTR_PT(882) <=
    Eq(( ROM_ADDR_L2(4) & ROM_ADDR_L2(5)
     ) , STD_ULOGIC_VECTOR'("00"));
MQQ1844:ROM32_INSTR_PT(883) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(5)
     ) , STD_ULOGIC_VECTOR'("00"));
MQQ1845:ROM32_INSTR_PT(884) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(5)
     ) , STD_ULOGIC_VECTOR'("0110"));
MQQ1846:ROM32_INSTR_PT(885) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) & ROM_ADDR_L2(5)
     ) , STD_ULOGIC_VECTOR'("0110"));
MQQ1847:ROM32_INSTR_PT(886) <=
    Eq(( ROM_ADDR_L2(3) & ROM_ADDR_L2(4) & 
    ROM_ADDR_L2(5) ) , STD_ULOGIC_VECTOR'("111"));
MQQ1848:ROM32_INSTR_PT(887) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(3) & 
    ROM_ADDR_L2(4) ) , STD_ULOGIC_VECTOR'("000"));
MQQ1849:ROM32_INSTR_PT(888) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(2) & 
    ROM_ADDR_L2(3) & ROM_ADDR_L2(4)
     ) , STD_ULOGIC_VECTOR'("0111"));
MQQ1850:ROM32_INSTR_PT(889) <=
    Eq(( ROM_ADDR_L2(0) & ROM_ADDR_L2(1) & 
    ROM_ADDR_L2(2) ) , STD_ULOGIC_VECTOR'("111"));
MQQ1851:ROM32_INSTR_PT(890) <=
    Eq(( ROM_ADDR_L2(2) ) , STD_ULOGIC'('1'));
MQQ1852:ROM32_INSTR_PT(891) <=
    Eq(( ROM_ADDR_L2(1) ) , STD_ULOGIC'('1'));
MQQ1853:ROM32_INSTR_PT(892) <=
    Eq(( ROM_ADDR_L2(0) ) , STD_ULOGIC'('0'));
MQQ1854:ROM32_INSTR_PT(893) <=
    '1';
MQQ1855:TEMPLATE(0) <= 
    (ROM32_INSTR_PT(28) OR ROM32_INSTR_PT(33)
     OR ROM32_INSTR_PT(45) OR ROM32_INSTR_PT(68)
     OR ROM32_INSTR_PT(76) OR ROM32_INSTR_PT(85)
     OR ROM32_INSTR_PT(113) OR ROM32_INSTR_PT(120)
     OR ROM32_INSTR_PT(128) OR ROM32_INSTR_PT(132)
     OR ROM32_INSTR_PT(142) OR ROM32_INSTR_PT(159)
     OR ROM32_INSTR_PT(162) OR ROM32_INSTR_PT(175)
     OR ROM32_INSTR_PT(176) OR ROM32_INSTR_PT(177)
     OR ROM32_INSTR_PT(180) OR ROM32_INSTR_PT(222)
     OR ROM32_INSTR_PT(226) OR ROM32_INSTR_PT(233)
     OR ROM32_INSTR_PT(237) OR ROM32_INSTR_PT(242)
     OR ROM32_INSTR_PT(255) OR ROM32_INSTR_PT(290)
     OR ROM32_INSTR_PT(292) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(335) OR ROM32_INSTR_PT(346)
     OR ROM32_INSTR_PT(351) OR ROM32_INSTR_PT(353)
     OR ROM32_INSTR_PT(356) OR ROM32_INSTR_PT(357)
     OR ROM32_INSTR_PT(359) OR ROM32_INSTR_PT(364)
     OR ROM32_INSTR_PT(365) OR ROM32_INSTR_PT(373)
     OR ROM32_INSTR_PT(381) OR ROM32_INSTR_PT(388)
     OR ROM32_INSTR_PT(391) OR ROM32_INSTR_PT(399)
     OR ROM32_INSTR_PT(425) OR ROM32_INSTR_PT(431)
     OR ROM32_INSTR_PT(467) OR ROM32_INSTR_PT(473)
     OR ROM32_INSTR_PT(527) OR ROM32_INSTR_PT(555)
     OR ROM32_INSTR_PT(563) OR ROM32_INSTR_PT(571)
     OR ROM32_INSTR_PT(586) OR ROM32_INSTR_PT(597)
     OR ROM32_INSTR_PT(604) OR ROM32_INSTR_PT(615)
     OR ROM32_INSTR_PT(652) OR ROM32_INSTR_PT(657)
     OR ROM32_INSTR_PT(664) OR ROM32_INSTR_PT(691)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(697)
     OR ROM32_INSTR_PT(711) OR ROM32_INSTR_PT(715)
     OR ROM32_INSTR_PT(716) OR ROM32_INSTR_PT(718)
     OR ROM32_INSTR_PT(729) OR ROM32_INSTR_PT(763)
     OR ROM32_INSTR_PT(792) OR ROM32_INSTR_PT(829)
     OR ROM32_INSTR_PT(831) OR ROM32_INSTR_PT(857)
     OR ROM32_INSTR_PT(872));
MQQ1856:TEMPLATE(1) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(7)
     OR ROM32_INSTR_PT(8) OR ROM32_INSTR_PT(9)
     OR ROM32_INSTR_PT(10) OR ROM32_INSTR_PT(13)
     OR ROM32_INSTR_PT(14) OR ROM32_INSTR_PT(16)
     OR ROM32_INSTR_PT(17) OR ROM32_INSTR_PT(20)
     OR ROM32_INSTR_PT(23) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(32) OR ROM32_INSTR_PT(35)
     OR ROM32_INSTR_PT(37) OR ROM32_INSTR_PT(39)
     OR ROM32_INSTR_PT(41) OR ROM32_INSTR_PT(42)
     OR ROM32_INSTR_PT(43) OR ROM32_INSTR_PT(49)
     OR ROM32_INSTR_PT(50) OR ROM32_INSTR_PT(51)
     OR ROM32_INSTR_PT(52) OR ROM32_INSTR_PT(53)
     OR ROM32_INSTR_PT(55) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(59)
     OR ROM32_INSTR_PT(63) OR ROM32_INSTR_PT(66)
     OR ROM32_INSTR_PT(67) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(73) OR ROM32_INSTR_PT(74)
     OR ROM32_INSTR_PT(77) OR ROM32_INSTR_PT(79)
     OR ROM32_INSTR_PT(80) OR ROM32_INSTR_PT(83)
     OR ROM32_INSTR_PT(84) OR ROM32_INSTR_PT(87)
     OR ROM32_INSTR_PT(90) OR ROM32_INSTR_PT(92)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(96)
     OR ROM32_INSTR_PT(97) OR ROM32_INSTR_PT(99)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(102) OR ROM32_INSTR_PT(103)
     OR ROM32_INSTR_PT(105) OR ROM32_INSTR_PT(106)
     OR ROM32_INSTR_PT(109) OR ROM32_INSTR_PT(110)
     OR ROM32_INSTR_PT(111) OR ROM32_INSTR_PT(114)
     OR ROM32_INSTR_PT(115) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(122) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(127) OR ROM32_INSTR_PT(130)
     OR ROM32_INSTR_PT(134) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(139) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(144) OR ROM32_INSTR_PT(148)
     OR ROM32_INSTR_PT(153) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(163) OR ROM32_INSTR_PT(164)
     OR ROM32_INSTR_PT(165) OR ROM32_INSTR_PT(169)
     OR ROM32_INSTR_PT(170) OR ROM32_INSTR_PT(171)
     OR ROM32_INSTR_PT(172) OR ROM32_INSTR_PT(179)
     OR ROM32_INSTR_PT(183) OR ROM32_INSTR_PT(184)
     OR ROM32_INSTR_PT(186) OR ROM32_INSTR_PT(192)
     OR ROM32_INSTR_PT(193) OR ROM32_INSTR_PT(195)
     OR ROM32_INSTR_PT(196) OR ROM32_INSTR_PT(199)
     OR ROM32_INSTR_PT(200) OR ROM32_INSTR_PT(202)
     OR ROM32_INSTR_PT(203) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(206) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(209) OR ROM32_INSTR_PT(215)
     OR ROM32_INSTR_PT(216) OR ROM32_INSTR_PT(218)
     OR ROM32_INSTR_PT(219) OR ROM32_INSTR_PT(220)
     OR ROM32_INSTR_PT(223) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(241)
     OR ROM32_INSTR_PT(243) OR ROM32_INSTR_PT(249)
     OR ROM32_INSTR_PT(250) OR ROM32_INSTR_PT(252)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(259)
     OR ROM32_INSTR_PT(260) OR ROM32_INSTR_PT(261)
     OR ROM32_INSTR_PT(262) OR ROM32_INSTR_PT(264)
     OR ROM32_INSTR_PT(267) OR ROM32_INSTR_PT(268)
     OR ROM32_INSTR_PT(269) OR ROM32_INSTR_PT(270)
     OR ROM32_INSTR_PT(273) OR ROM32_INSTR_PT(274)
     OR ROM32_INSTR_PT(275) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(280) OR ROM32_INSTR_PT(282)
     OR ROM32_INSTR_PT(283) OR ROM32_INSTR_PT(284)
     OR ROM32_INSTR_PT(287) OR ROM32_INSTR_PT(288)
     OR ROM32_INSTR_PT(289) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(306) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(321) OR ROM32_INSTR_PT(323)
     OR ROM32_INSTR_PT(328) OR ROM32_INSTR_PT(331)
     OR ROM32_INSTR_PT(342) OR ROM32_INSTR_PT(345)
     OR ROM32_INSTR_PT(348) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(352) OR ROM32_INSTR_PT(355)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(362)
     OR ROM32_INSTR_PT(363) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(368)
     OR ROM32_INSTR_PT(370) OR ROM32_INSTR_PT(371)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(382)
     OR ROM32_INSTR_PT(383) OR ROM32_INSTR_PT(386)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(390)
     OR ROM32_INSTR_PT(392) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(396) OR ROM32_INSTR_PT(400)
     OR ROM32_INSTR_PT(401) OR ROM32_INSTR_PT(402)
     OR ROM32_INSTR_PT(404) OR ROM32_INSTR_PT(405)
     OR ROM32_INSTR_PT(406) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(411) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(417)
     OR ROM32_INSTR_PT(418) OR ROM32_INSTR_PT(421)
     OR ROM32_INSTR_PT(422) OR ROM32_INSTR_PT(423)
     OR ROM32_INSTR_PT(424) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(428) OR ROM32_INSTR_PT(430)
     OR ROM32_INSTR_PT(433) OR ROM32_INSTR_PT(434)
     OR ROM32_INSTR_PT(435) OR ROM32_INSTR_PT(436)
     OR ROM32_INSTR_PT(438) OR ROM32_INSTR_PT(441)
     OR ROM32_INSTR_PT(442) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(452)
     OR ROM32_INSTR_PT(453) OR ROM32_INSTR_PT(454)
     OR ROM32_INSTR_PT(458) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(464) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(474)
     OR ROM32_INSTR_PT(475) OR ROM32_INSTR_PT(476)
     OR ROM32_INSTR_PT(477) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(480)
     OR ROM32_INSTR_PT(481) OR ROM32_INSTR_PT(482)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(491) OR ROM32_INSTR_PT(494)
     OR ROM32_INSTR_PT(496) OR ROM32_INSTR_PT(497)
     OR ROM32_INSTR_PT(498) OR ROM32_INSTR_PT(501)
     OR ROM32_INSTR_PT(502) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(505) OR ROM32_INSTR_PT(506)
     OR ROM32_INSTR_PT(507) OR ROM32_INSTR_PT(508)
     OR ROM32_INSTR_PT(509) OR ROM32_INSTR_PT(514)
     OR ROM32_INSTR_PT(517) OR ROM32_INSTR_PT(519)
     OR ROM32_INSTR_PT(520) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(524)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(531)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(535) OR ROM32_INSTR_PT(536)
     OR ROM32_INSTR_PT(538) OR ROM32_INSTR_PT(539)
     OR ROM32_INSTR_PT(541) OR ROM32_INSTR_PT(543)
     OR ROM32_INSTR_PT(544) OR ROM32_INSTR_PT(546)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(550)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(556)
     OR ROM32_INSTR_PT(557) OR ROM32_INSTR_PT(558)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(566)
     OR ROM32_INSTR_PT(568) OR ROM32_INSTR_PT(569)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(575) OR ROM32_INSTR_PT(578)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(580)
     OR ROM32_INSTR_PT(581) OR ROM32_INSTR_PT(582)
     OR ROM32_INSTR_PT(583) OR ROM32_INSTR_PT(584)
     OR ROM32_INSTR_PT(585) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(589) OR ROM32_INSTR_PT(590)
     OR ROM32_INSTR_PT(593) OR ROM32_INSTR_PT(595)
     OR ROM32_INSTR_PT(598) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(601)
     OR ROM32_INSTR_PT(602) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(606) OR ROM32_INSTR_PT(607)
     OR ROM32_INSTR_PT(608) OR ROM32_INSTR_PT(609)
     OR ROM32_INSTR_PT(610) OR ROM32_INSTR_PT(611)
     OR ROM32_INSTR_PT(612) OR ROM32_INSTR_PT(613)
     OR ROM32_INSTR_PT(614) OR ROM32_INSTR_PT(620)
     OR ROM32_INSTR_PT(621) OR ROM32_INSTR_PT(624)
     OR ROM32_INSTR_PT(625) OR ROM32_INSTR_PT(626)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(634)
     OR ROM32_INSTR_PT(635) OR ROM32_INSTR_PT(638)
     OR ROM32_INSTR_PT(639) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(643) OR ROM32_INSTR_PT(644)
     OR ROM32_INSTR_PT(647) OR ROM32_INSTR_PT(654)
     OR ROM32_INSTR_PT(660) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(666) OR ROM32_INSTR_PT(674)
     OR ROM32_INSTR_PT(677) OR ROM32_INSTR_PT(678)
     OR ROM32_INSTR_PT(680) OR ROM32_INSTR_PT(684)
     OR ROM32_INSTR_PT(685) OR ROM32_INSTR_PT(698)
     OR ROM32_INSTR_PT(708) OR ROM32_INSTR_PT(713)
     OR ROM32_INSTR_PT(719) OR ROM32_INSTR_PT(726)
     OR ROM32_INSTR_PT(733) OR ROM32_INSTR_PT(736)
     OR ROM32_INSTR_PT(745) OR ROM32_INSTR_PT(755)
     OR ROM32_INSTR_PT(762) OR ROM32_INSTR_PT(770)
     OR ROM32_INSTR_PT(785) OR ROM32_INSTR_PT(795)
     OR ROM32_INSTR_PT(801) OR ROM32_INSTR_PT(805)
     OR ROM32_INSTR_PT(812) OR ROM32_INSTR_PT(817)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(845)
     OR ROM32_INSTR_PT(847) OR ROM32_INSTR_PT(851)
     OR ROM32_INSTR_PT(853) OR ROM32_INSTR_PT(854)
     OR ROM32_INSTR_PT(855) OR ROM32_INSTR_PT(862)
     OR ROM32_INSTR_PT(869) OR ROM32_INSTR_PT(870)
     OR ROM32_INSTR_PT(871) OR ROM32_INSTR_PT(878)
     OR ROM32_INSTR_PT(889));
MQQ1857:TEMPLATE(2) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(7)
     OR ROM32_INSTR_PT(13) OR ROM32_INSTR_PT(14)
     OR ROM32_INSTR_PT(18) OR ROM32_INSTR_PT(23)
     OR ROM32_INSTR_PT(27) OR ROM32_INSTR_PT(29)
     OR ROM32_INSTR_PT(31) OR ROM32_INSTR_PT(35)
     OR ROM32_INSTR_PT(38) OR ROM32_INSTR_PT(39)
     OR ROM32_INSTR_PT(41) OR ROM32_INSTR_PT(42)
     OR ROM32_INSTR_PT(43) OR ROM32_INSTR_PT(53)
     OR ROM32_INSTR_PT(56) OR ROM32_INSTR_PT(57)
     OR ROM32_INSTR_PT(62) OR ROM32_INSTR_PT(70)
     OR ROM32_INSTR_PT(72) OR ROM32_INSTR_PT(79)
     OR ROM32_INSTR_PT(80) OR ROM32_INSTR_PT(81)
     OR ROM32_INSTR_PT(83) OR ROM32_INSTR_PT(92)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(98) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(102) OR ROM32_INSTR_PT(105)
     OR ROM32_INSTR_PT(109) OR ROM32_INSTR_PT(110)
     OR ROM32_INSTR_PT(111) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(122) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(130) OR ROM32_INSTR_PT(139)
     OR ROM32_INSTR_PT(141) OR ROM32_INSTR_PT(144)
     OR ROM32_INSTR_PT(145) OR ROM32_INSTR_PT(146)
     OR ROM32_INSTR_PT(147) OR ROM32_INSTR_PT(150)
     OR ROM32_INSTR_PT(151) OR ROM32_INSTR_PT(153)
     OR ROM32_INSTR_PT(158) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(165) OR ROM32_INSTR_PT(166)
     OR ROM32_INSTR_PT(172) OR ROM32_INSTR_PT(174)
     OR ROM32_INSTR_PT(185) OR ROM32_INSTR_PT(186)
     OR ROM32_INSTR_PT(187) OR ROM32_INSTR_PT(189)
     OR ROM32_INSTR_PT(192) OR ROM32_INSTR_PT(193)
     OR ROM32_INSTR_PT(195) OR ROM32_INSTR_PT(199)
     OR ROM32_INSTR_PT(203) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(206) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(208) OR ROM32_INSTR_PT(209)
     OR ROM32_INSTR_PT(210) OR ROM32_INSTR_PT(218)
     OR ROM32_INSTR_PT(228) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(230) OR ROM32_INSTR_PT(232)
     OR ROM32_INSTR_PT(235) OR ROM32_INSTR_PT(240)
     OR ROM32_INSTR_PT(245) OR ROM32_INSTR_PT(249)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(252)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(262)
     OR ROM32_INSTR_PT(268) OR ROM32_INSTR_PT(275)
     OR ROM32_INSTR_PT(279) OR ROM32_INSTR_PT(285)
     OR ROM32_INSTR_PT(287) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(291) OR ROM32_INSTR_PT(294)
     OR ROM32_INSTR_PT(302) OR ROM32_INSTR_PT(305)
     OR ROM32_INSTR_PT(307) OR ROM32_INSTR_PT(311)
     OR ROM32_INSTR_PT(322) OR ROM32_INSTR_PT(323)
     OR ROM32_INSTR_PT(325) OR ROM32_INSTR_PT(329)
     OR ROM32_INSTR_PT(331) OR ROM32_INSTR_PT(332)
     OR ROM32_INSTR_PT(337) OR ROM32_INSTR_PT(338)
     OR ROM32_INSTR_PT(339) OR ROM32_INSTR_PT(342)
     OR ROM32_INSTR_PT(350) OR ROM32_INSTR_PT(352)
     OR ROM32_INSTR_PT(355) OR ROM32_INSTR_PT(362)
     OR ROM32_INSTR_PT(363) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(368)
     OR ROM32_INSTR_PT(370) OR ROM32_INSTR_PT(374)
     OR ROM32_INSTR_PT(376) OR ROM32_INSTR_PT(378)
     OR ROM32_INSTR_PT(382) OR ROM32_INSTR_PT(386)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(393)
     OR ROM32_INSTR_PT(394) OR ROM32_INSTR_PT(395)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(400)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(404)
     OR ROM32_INSTR_PT(405) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(416)
     OR ROM32_INSTR_PT(417) OR ROM32_INSTR_PT(418)
     OR ROM32_INSTR_PT(419) OR ROM32_INSTR_PT(422)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(435)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(438)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(442)
     OR ROM32_INSTR_PT(443) OR ROM32_INSTR_PT(446)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(452)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(456)
     OR ROM32_INSTR_PT(458) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(463) OR ROM32_INSTR_PT(464)
     OR ROM32_INSTR_PT(465) OR ROM32_INSTR_PT(468)
     OR ROM32_INSTR_PT(469) OR ROM32_INSTR_PT(471)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(474)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(480)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(489)
     OR ROM32_INSTR_PT(496) OR ROM32_INSTR_PT(497)
     OR ROM32_INSTR_PT(498) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(505) OR ROM32_INSTR_PT(507)
     OR ROM32_INSTR_PT(513) OR ROM32_INSTR_PT(514)
     OR ROM32_INSTR_PT(517) OR ROM32_INSTR_PT(532)
     OR ROM32_INSTR_PT(537) OR ROM32_INSTR_PT(539)
     OR ROM32_INSTR_PT(541) OR ROM32_INSTR_PT(544)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(549)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(561)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(569)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(577) OR ROM32_INSTR_PT(579)
     OR ROM32_INSTR_PT(580) OR ROM32_INSTR_PT(584)
     OR ROM32_INSTR_PT(587) OR ROM32_INSTR_PT(589)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(593)
     OR ROM32_INSTR_PT(596) OR ROM32_INSTR_PT(598)
     OR ROM32_INSTR_PT(599) OR ROM32_INSTR_PT(600)
     OR ROM32_INSTR_PT(605) OR ROM32_INSTR_PT(606)
     OR ROM32_INSTR_PT(607) OR ROM32_INSTR_PT(608)
     OR ROM32_INSTR_PT(609) OR ROM32_INSTR_PT(610)
     OR ROM32_INSTR_PT(611) OR ROM32_INSTR_PT(614)
     OR ROM32_INSTR_PT(620) OR ROM32_INSTR_PT(624)
     OR ROM32_INSTR_PT(625) OR ROM32_INSTR_PT(629)
     OR ROM32_INSTR_PT(632) OR ROM32_INSTR_PT(634)
     OR ROM32_INSTR_PT(638) OR ROM32_INSTR_PT(640)
     OR ROM32_INSTR_PT(643) OR ROM32_INSTR_PT(653)
     OR ROM32_INSTR_PT(659) OR ROM32_INSTR_PT(660)
     OR ROM32_INSTR_PT(663) OR ROM32_INSTR_PT(668)
     OR ROM32_INSTR_PT(672) OR ROM32_INSTR_PT(678)
     OR ROM32_INSTR_PT(680) OR ROM32_INSTR_PT(684)
     OR ROM32_INSTR_PT(685) OR ROM32_INSTR_PT(689)
     OR ROM32_INSTR_PT(698) OR ROM32_INSTR_PT(704)
     OR ROM32_INSTR_PT(705) OR ROM32_INSTR_PT(708)
     OR ROM32_INSTR_PT(713) OR ROM32_INSTR_PT(720)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(733)
     OR ROM32_INSTR_PT(751) OR ROM32_INSTR_PT(752)
     OR ROM32_INSTR_PT(753) OR ROM32_INSTR_PT(759)
     OR ROM32_INSTR_PT(774) OR ROM32_INSTR_PT(785)
     OR ROM32_INSTR_PT(787) OR ROM32_INSTR_PT(790)
     OR ROM32_INSTR_PT(795) OR ROM32_INSTR_PT(799)
     OR ROM32_INSTR_PT(801) OR ROM32_INSTR_PT(803)
     OR ROM32_INSTR_PT(805) OR ROM32_INSTR_PT(807)
     OR ROM32_INSTR_PT(812) OR ROM32_INSTR_PT(817)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(823)
     OR ROM32_INSTR_PT(845) OR ROM32_INSTR_PT(847)
     OR ROM32_INSTR_PT(851) OR ROM32_INSTR_PT(853)
     OR ROM32_INSTR_PT(854) OR ROM32_INSTR_PT(869)
     OR ROM32_INSTR_PT(871) OR ROM32_INSTR_PT(878)
     OR ROM32_INSTR_PT(881) OR ROM32_INSTR_PT(889)
    );
MQQ1858:TEMPLATE(3) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(7)
     OR ROM32_INSTR_PT(8) OR ROM32_INSTR_PT(9)
     OR ROM32_INSTR_PT(10) OR ROM32_INSTR_PT(13)
     OR ROM32_INSTR_PT(14) OR ROM32_INSTR_PT(16)
     OR ROM32_INSTR_PT(17) OR ROM32_INSTR_PT(18)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(23)
     OR ROM32_INSTR_PT(26) OR ROM32_INSTR_PT(27)
     OR ROM32_INSTR_PT(28) OR ROM32_INSTR_PT(31)
     OR ROM32_INSTR_PT(32) OR ROM32_INSTR_PT(33)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(37)
     OR ROM32_INSTR_PT(38) OR ROM32_INSTR_PT(39)
     OR ROM32_INSTR_PT(41) OR ROM32_INSTR_PT(42)
     OR ROM32_INSTR_PT(43) OR ROM32_INSTR_PT(45)
     OR ROM32_INSTR_PT(49) OR ROM32_INSTR_PT(52)
     OR ROM32_INSTR_PT(53) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(59)
     OR ROM32_INSTR_PT(62) OR ROM32_INSTR_PT(63)
     OR ROM32_INSTR_PT(66) OR ROM32_INSTR_PT(67)
     OR ROM32_INSTR_PT(70) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(73) OR ROM32_INSTR_PT(74)
     OR ROM32_INSTR_PT(77) OR ROM32_INSTR_PT(78)
     OR ROM32_INSTR_PT(79) OR ROM32_INSTR_PT(80)
     OR ROM32_INSTR_PT(83) OR ROM32_INSTR_PT(84)
     OR ROM32_INSTR_PT(85) OR ROM32_INSTR_PT(87)
     OR ROM32_INSTR_PT(90) OR ROM32_INSTR_PT(92)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(97) OR ROM32_INSTR_PT(98)
     OR ROM32_INSTR_PT(99) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(102) OR ROM32_INSTR_PT(103)
     OR ROM32_INSTR_PT(105) OR ROM32_INSTR_PT(109)
     OR ROM32_INSTR_PT(110) OR ROM32_INSTR_PT(111)
     OR ROM32_INSTR_PT(114) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(122) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(127) OR ROM32_INSTR_PT(130)
     OR ROM32_INSTR_PT(131) OR ROM32_INSTR_PT(134)
     OR ROM32_INSTR_PT(139) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(144) OR ROM32_INSTR_PT(145)
     OR ROM32_INSTR_PT(146) OR ROM32_INSTR_PT(147)
     OR ROM32_INSTR_PT(148) OR ROM32_INSTR_PT(150)
     OR ROM32_INSTR_PT(151) OR ROM32_INSTR_PT(153)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(162) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(164) OR ROM32_INSTR_PT(165)
     OR ROM32_INSTR_PT(166) OR ROM32_INSTR_PT(169)
     OR ROM32_INSTR_PT(171) OR ROM32_INSTR_PT(172)
     OR ROM32_INSTR_PT(173) OR ROM32_INSTR_PT(174)
     OR ROM32_INSTR_PT(176) OR ROM32_INSTR_PT(177)
     OR ROM32_INSTR_PT(178) OR ROM32_INSTR_PT(179)
     OR ROM32_INSTR_PT(180) OR ROM32_INSTR_PT(181)
     OR ROM32_INSTR_PT(184) OR ROM32_INSTR_PT(185)
     OR ROM32_INSTR_PT(186) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(189) OR ROM32_INSTR_PT(192)
     OR ROM32_INSTR_PT(194) OR ROM32_INSTR_PT(199)
     OR ROM32_INSTR_PT(200) OR ROM32_INSTR_PT(202)
     OR ROM32_INSTR_PT(203) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(206) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(208) OR ROM32_INSTR_PT(209)
     OR ROM32_INSTR_PT(210) OR ROM32_INSTR_PT(212)
     OR ROM32_INSTR_PT(216) OR ROM32_INSTR_PT(218)
     OR ROM32_INSTR_PT(219) OR ROM32_INSTR_PT(220)
     OR ROM32_INSTR_PT(222) OR ROM32_INSTR_PT(223)
     OR ROM32_INSTR_PT(224) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(228)
     OR ROM32_INSTR_PT(229) OR ROM32_INSTR_PT(230)
     OR ROM32_INSTR_PT(232) OR ROM32_INSTR_PT(233)
     OR ROM32_INSTR_PT(235) OR ROM32_INSTR_PT(238)
     OR ROM32_INSTR_PT(240) OR ROM32_INSTR_PT(242)
     OR ROM32_INSTR_PT(244) OR ROM32_INSTR_PT(245)
     OR ROM32_INSTR_PT(249) OR ROM32_INSTR_PT(250)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(252)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(255)
     OR ROM32_INSTR_PT(256) OR ROM32_INSTR_PT(257)
     OR ROM32_INSTR_PT(259) OR ROM32_INSTR_PT(261)
     OR ROM32_INSTR_PT(262) OR ROM32_INSTR_PT(264)
     OR ROM32_INSTR_PT(266) OR ROM32_INSTR_PT(267)
     OR ROM32_INSTR_PT(268) OR ROM32_INSTR_PT(269)
     OR ROM32_INSTR_PT(270) OR ROM32_INSTR_PT(271)
     OR ROM32_INSTR_PT(272) OR ROM32_INSTR_PT(273)
     OR ROM32_INSTR_PT(275) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(279) OR ROM32_INSTR_PT(280)
     OR ROM32_INSTR_PT(284) OR ROM32_INSTR_PT(285)
     OR ROM32_INSTR_PT(288) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(290) OR ROM32_INSTR_PT(291)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(302)
     OR ROM32_INSTR_PT(303) OR ROM32_INSTR_PT(305)
     OR ROM32_INSTR_PT(307) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(311) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(322)
     OR ROM32_INSTR_PT(323) OR ROM32_INSTR_PT(325)
     OR ROM32_INSTR_PT(328) OR ROM32_INSTR_PT(329)
     OR ROM32_INSTR_PT(332) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(337) OR ROM32_INSTR_PT(338)
     OR ROM32_INSTR_PT(339) OR ROM32_INSTR_PT(344)
     OR ROM32_INSTR_PT(346) OR ROM32_INSTR_PT(348)
     OR ROM32_INSTR_PT(350) OR ROM32_INSTR_PT(357)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(362)
     OR ROM32_INSTR_PT(363) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(368)
     OR ROM32_INSTR_PT(371) OR ROM32_INSTR_PT(373)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(378) OR ROM32_INSTR_PT(379)
     OR ROM32_INSTR_PT(381) OR ROM32_INSTR_PT(382)
     OR ROM32_INSTR_PT(383) OR ROM32_INSTR_PT(386)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(388)
     OR ROM32_INSTR_PT(390) OR ROM32_INSTR_PT(392)
     OR ROM32_INSTR_PT(393) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(395) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(400)
     OR ROM32_INSTR_PT(401) OR ROM32_INSTR_PT(402)
     OR ROM32_INSTR_PT(404) OR ROM32_INSTR_PT(405)
     OR ROM32_INSTR_PT(406) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(411) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(416)
     OR ROM32_INSTR_PT(417) OR ROM32_INSTR_PT(418)
     OR ROM32_INSTR_PT(419) OR ROM32_INSTR_PT(421)
     OR ROM32_INSTR_PT(422) OR ROM32_INSTR_PT(423)
     OR ROM32_INSTR_PT(424) OR ROM32_INSTR_PT(425)
     OR ROM32_INSTR_PT(426) OR ROM32_INSTR_PT(433)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(435)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(437)
     OR ROM32_INSTR_PT(438) OR ROM32_INSTR_PT(441)
     OR ROM32_INSTR_PT(442) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(446) OR ROM32_INSTR_PT(451)
     OR ROM32_INSTR_PT(452) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(456)
     OR ROM32_INSTR_PT(458) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(463) OR ROM32_INSTR_PT(464)
     OR ROM32_INSTR_PT(465) OR ROM32_INSTR_PT(467)
     OR ROM32_INSTR_PT(468) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(471) OR ROM32_INSTR_PT(472)
     OR ROM32_INSTR_PT(474) OR ROM32_INSTR_PT(475)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(480)
     OR ROM32_INSTR_PT(481) OR ROM32_INSTR_PT(482)
     OR ROM32_INSTR_PT(484) OR ROM32_INSTR_PT(486)
     OR ROM32_INSTR_PT(489) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(494) OR ROM32_INSTR_PT(495)
     OR ROM32_INSTR_PT(496) OR ROM32_INSTR_PT(497)
     OR ROM32_INSTR_PT(502) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(505) OR ROM32_INSTR_PT(506)
     OR ROM32_INSTR_PT(507) OR ROM32_INSTR_PT(508)
     OR ROM32_INSTR_PT(513) OR ROM32_INSTR_PT(514)
     OR ROM32_INSTR_PT(517) OR ROM32_INSTR_PT(519)
     OR ROM32_INSTR_PT(520) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(524)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(537) OR ROM32_INSTR_PT(539)
     OR ROM32_INSTR_PT(541) OR ROM32_INSTR_PT(544)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(549)
     OR ROM32_INSTR_PT(550) OR ROM32_INSTR_PT(551)
     OR ROM32_INSTR_PT(552) OR ROM32_INSTR_PT(554)
     OR ROM32_INSTR_PT(556) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(561)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(568)
     OR ROM32_INSTR_PT(569) OR ROM32_INSTR_PT(570)
     OR ROM32_INSTR_PT(571) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(575) OR ROM32_INSTR_PT(577)
     OR ROM32_INSTR_PT(578) OR ROM32_INSTR_PT(579)
     OR ROM32_INSTR_PT(580) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(582) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(584) OR ROM32_INSTR_PT(585)
     OR ROM32_INSTR_PT(586) OR ROM32_INSTR_PT(587)
     OR ROM32_INSTR_PT(588) OR ROM32_INSTR_PT(590)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(593)
     OR ROM32_INSTR_PT(595) OR ROM32_INSTR_PT(596)
     OR ROM32_INSTR_PT(598) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(602)
     OR ROM32_INSTR_PT(604) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(606) OR ROM32_INSTR_PT(607)
     OR ROM32_INSTR_PT(608) OR ROM32_INSTR_PT(609)
     OR ROM32_INSTR_PT(610) OR ROM32_INSTR_PT(611)
     OR ROM32_INSTR_PT(612) OR ROM32_INSTR_PT(614)
     OR ROM32_INSTR_PT(620) OR ROM32_INSTR_PT(621)
     OR ROM32_INSTR_PT(624) OR ROM32_INSTR_PT(625)
     OR ROM32_INSTR_PT(626) OR ROM32_INSTR_PT(629)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(632)
     OR ROM32_INSTR_PT(634) OR ROM32_INSTR_PT(638)
     OR ROM32_INSTR_PT(639) OR ROM32_INSTR_PT(640)
     OR ROM32_INSTR_PT(642) OR ROM32_INSTR_PT(643)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(653)
     OR ROM32_INSTR_PT(657) OR ROM32_INSTR_PT(659)
     OR ROM32_INSTR_PT(660) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(664) OR ROM32_INSTR_PT(666)
     OR ROM32_INSTR_PT(668) OR ROM32_INSTR_PT(672)
     OR ROM32_INSTR_PT(677) OR ROM32_INSTR_PT(680)
     OR ROM32_INSTR_PT(684) OR ROM32_INSTR_PT(689)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(698)
     OR ROM32_INSTR_PT(702) OR ROM32_INSTR_PT(704)
     OR ROM32_INSTR_PT(708) OR ROM32_INSTR_PT(713)
     OR ROM32_INSTR_PT(718) OR ROM32_INSTR_PT(719)
     OR ROM32_INSTR_PT(720) OR ROM32_INSTR_PT(726)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(729)
     OR ROM32_INSTR_PT(736) OR ROM32_INSTR_PT(751)
     OR ROM32_INSTR_PT(752) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(755) OR ROM32_INSTR_PT(759)
     OR ROM32_INSTR_PT(762) OR ROM32_INSTR_PT(770)
     OR ROM32_INSTR_PT(774) OR ROM32_INSTR_PT(787)
     OR ROM32_INSTR_PT(790) OR ROM32_INSTR_PT(792)
     OR ROM32_INSTR_PT(803) OR ROM32_INSTR_PT(805)
     OR ROM32_INSTR_PT(807) OR ROM32_INSTR_PT(812)
     OR ROM32_INSTR_PT(817) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(823) OR ROM32_INSTR_PT(831)
     OR ROM32_INSTR_PT(845) OR ROM32_INSTR_PT(853)
     OR ROM32_INSTR_PT(854) OR ROM32_INSTR_PT(855)
     OR ROM32_INSTR_PT(857) OR ROM32_INSTR_PT(862)
     OR ROM32_INSTR_PT(869) OR ROM32_INSTR_PT(870)
     OR ROM32_INSTR_PT(878) OR ROM32_INSTR_PT(881)
    );
MQQ1859:TEMPLATE(4) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(7)
     OR ROM32_INSTR_PT(13) OR ROM32_INSTR_PT(14)
     OR ROM32_INSTR_PT(18) OR ROM32_INSTR_PT(23)
     OR ROM32_INSTR_PT(27) OR ROM32_INSTR_PT(28)
     OR ROM32_INSTR_PT(29) OR ROM32_INSTR_PT(31)
     OR ROM32_INSTR_PT(33) OR ROM32_INSTR_PT(35)
     OR ROM32_INSTR_PT(38) OR ROM32_INSTR_PT(39)
     OR ROM32_INSTR_PT(41) OR ROM32_INSTR_PT(42)
     OR ROM32_INSTR_PT(43) OR ROM32_INSTR_PT(45)
     OR ROM32_INSTR_PT(53) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(62)
     OR ROM32_INSTR_PT(68) OR ROM32_INSTR_PT(70)
     OR ROM32_INSTR_PT(72) OR ROM32_INSTR_PT(76)
     OR ROM32_INSTR_PT(79) OR ROM32_INSTR_PT(80)
     OR ROM32_INSTR_PT(81) OR ROM32_INSTR_PT(83)
     OR ROM32_INSTR_PT(85) OR ROM32_INSTR_PT(92)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(98) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(102) OR ROM32_INSTR_PT(105)
     OR ROM32_INSTR_PT(109) OR ROM32_INSTR_PT(110)
     OR ROM32_INSTR_PT(111) OR ROM32_INSTR_PT(113)
     OR ROM32_INSTR_PT(117) OR ROM32_INSTR_PT(120)
     OR ROM32_INSTR_PT(122) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(128) OR ROM32_INSTR_PT(130)
     OR ROM32_INSTR_PT(138) OR ROM32_INSTR_PT(139)
     OR ROM32_INSTR_PT(141) OR ROM32_INSTR_PT(142)
     OR ROM32_INSTR_PT(144) OR ROM32_INSTR_PT(145)
     OR ROM32_INSTR_PT(146) OR ROM32_INSTR_PT(147)
     OR ROM32_INSTR_PT(150) OR ROM32_INSTR_PT(151)
     OR ROM32_INSTR_PT(153) OR ROM32_INSTR_PT(155)
     OR ROM32_INSTR_PT(158) OR ROM32_INSTR_PT(159)
     OR ROM32_INSTR_PT(162) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(165) OR ROM32_INSTR_PT(166)
     OR ROM32_INSTR_PT(172) OR ROM32_INSTR_PT(173)
     OR ROM32_INSTR_PT(174) OR ROM32_INSTR_PT(175)
     OR ROM32_INSTR_PT(176) OR ROM32_INSTR_PT(177)
     OR ROM32_INSTR_PT(178) OR ROM32_INSTR_PT(180)
     OR ROM32_INSTR_PT(181) OR ROM32_INSTR_PT(185)
     OR ROM32_INSTR_PT(186) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(189) OR ROM32_INSTR_PT(192)
     OR ROM32_INSTR_PT(193) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(199) OR ROM32_INSTR_PT(203)
     OR ROM32_INSTR_PT(205) OR ROM32_INSTR_PT(206)
     OR ROM32_INSTR_PT(207) OR ROM32_INSTR_PT(208)
     OR ROM32_INSTR_PT(209) OR ROM32_INSTR_PT(210)
     OR ROM32_INSTR_PT(212) OR ROM32_INSTR_PT(218)
     OR ROM32_INSTR_PT(222) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(228) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(230) OR ROM32_INSTR_PT(232)
     OR ROM32_INSTR_PT(233) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(237) OR ROM32_INSTR_PT(240)
     OR ROM32_INSTR_PT(242) OR ROM32_INSTR_PT(245)
     OR ROM32_INSTR_PT(249) OR ROM32_INSTR_PT(251)
     OR ROM32_INSTR_PT(252) OR ROM32_INSTR_PT(254)
     OR ROM32_INSTR_PT(255) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(262)
     OR ROM32_INSTR_PT(266) OR ROM32_INSTR_PT(268)
     OR ROM32_INSTR_PT(272) OR ROM32_INSTR_PT(275)
     OR ROM32_INSTR_PT(279) OR ROM32_INSTR_PT(285)
     OR ROM32_INSTR_PT(287) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(290) OR ROM32_INSTR_PT(291)
     OR ROM32_INSTR_PT(292) OR ROM32_INSTR_PT(294)
     OR ROM32_INSTR_PT(302) OR ROM32_INSTR_PT(305)
     OR ROM32_INSTR_PT(307) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(311) OR ROM32_INSTR_PT(318)
     OR ROM32_INSTR_PT(322) OR ROM32_INSTR_PT(323)
     OR ROM32_INSTR_PT(325) OR ROM32_INSTR_PT(329)
     OR ROM32_INSTR_PT(332) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(337) OR ROM32_INSTR_PT(338)
     OR ROM32_INSTR_PT(339) OR ROM32_INSTR_PT(344)
     OR ROM32_INSTR_PT(346) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(356) OR ROM32_INSTR_PT(357)
     OR ROM32_INSTR_PT(358) OR ROM32_INSTR_PT(359)
     OR ROM32_INSTR_PT(362) OR ROM32_INSTR_PT(363)
     OR ROM32_INSTR_PT(365) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(368)
     OR ROM32_INSTR_PT(370) OR ROM32_INSTR_PT(373)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(378) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(382) OR ROM32_INSTR_PT(386)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(388)
     OR ROM32_INSTR_PT(391) OR ROM32_INSTR_PT(393)
     OR ROM32_INSTR_PT(394) OR ROM32_INSTR_PT(395)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(399)
     OR ROM32_INSTR_PT(400) OR ROM32_INSTR_PT(402)
     OR ROM32_INSTR_PT(404) OR ROM32_INSTR_PT(405)
     OR ROM32_INSTR_PT(409) OR ROM32_INSTR_PT(415)
     OR ROM32_INSTR_PT(416) OR ROM32_INSTR_PT(417)
     OR ROM32_INSTR_PT(418) OR ROM32_INSTR_PT(419)
     OR ROM32_INSTR_PT(422) OR ROM32_INSTR_PT(423)
     OR ROM32_INSTR_PT(425) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(435)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(438)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(442)
     OR ROM32_INSTR_PT(443) OR ROM32_INSTR_PT(446)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(452)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(456)
     OR ROM32_INSTR_PT(458) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(463) OR ROM32_INSTR_PT(464)
     OR ROM32_INSTR_PT(465) OR ROM32_INSTR_PT(467)
     OR ROM32_INSTR_PT(468) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(471) OR ROM32_INSTR_PT(472)
     OR ROM32_INSTR_PT(473) OR ROM32_INSTR_PT(474)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(480)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(489)
     OR ROM32_INSTR_PT(496) OR ROM32_INSTR_PT(497)
     OR ROM32_INSTR_PT(498) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(505) OR ROM32_INSTR_PT(507)
     OR ROM32_INSTR_PT(513) OR ROM32_INSTR_PT(514)
     OR ROM32_INSTR_PT(517) OR ROM32_INSTR_PT(527)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(537)
     OR ROM32_INSTR_PT(539) OR ROM32_INSTR_PT(541)
     OR ROM32_INSTR_PT(544) OR ROM32_INSTR_PT(547)
     OR ROM32_INSTR_PT(549) OR ROM32_INSTR_PT(551)
     OR ROM32_INSTR_PT(555) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(561)
     OR ROM32_INSTR_PT(563) OR ROM32_INSTR_PT(566)
     OR ROM32_INSTR_PT(569) OR ROM32_INSTR_PT(570)
     OR ROM32_INSTR_PT(571) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(577) OR ROM32_INSTR_PT(579)
     OR ROM32_INSTR_PT(580) OR ROM32_INSTR_PT(584)
     OR ROM32_INSTR_PT(586) OR ROM32_INSTR_PT(587)
     OR ROM32_INSTR_PT(589) OR ROM32_INSTR_PT(591)
     OR ROM32_INSTR_PT(593) OR ROM32_INSTR_PT(596)
     OR ROM32_INSTR_PT(597) OR ROM32_INSTR_PT(598)
     OR ROM32_INSTR_PT(599) OR ROM32_INSTR_PT(600)
     OR ROM32_INSTR_PT(604) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(606) OR ROM32_INSTR_PT(607)
     OR ROM32_INSTR_PT(608) OR ROM32_INSTR_PT(609)
     OR ROM32_INSTR_PT(610) OR ROM32_INSTR_PT(611)
     OR ROM32_INSTR_PT(614) OR ROM32_INSTR_PT(620)
     OR ROM32_INSTR_PT(624) OR ROM32_INSTR_PT(625)
     OR ROM32_INSTR_PT(629) OR ROM32_INSTR_PT(632)
     OR ROM32_INSTR_PT(634) OR ROM32_INSTR_PT(638)
     OR ROM32_INSTR_PT(640) OR ROM32_INSTR_PT(641)
     OR ROM32_INSTR_PT(643) OR ROM32_INSTR_PT(652)
     OR ROM32_INSTR_PT(653) OR ROM32_INSTR_PT(659)
     OR ROM32_INSTR_PT(660) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(664) OR ROM32_INSTR_PT(668)
     OR ROM32_INSTR_PT(672) OR ROM32_INSTR_PT(680)
     OR ROM32_INSTR_PT(683) OR ROM32_INSTR_PT(684)
     OR ROM32_INSTR_PT(689) OR ROM32_INSTR_PT(691)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(697)
     OR ROM32_INSTR_PT(698) OR ROM32_INSTR_PT(702)
     OR ROM32_INSTR_PT(704) OR ROM32_INSTR_PT(708)
     OR ROM32_INSTR_PT(711) OR ROM32_INSTR_PT(713)
     OR ROM32_INSTR_PT(718) OR ROM32_INSTR_PT(720)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(729)
     OR ROM32_INSTR_PT(733) OR ROM32_INSTR_PT(751)
     OR ROM32_INSTR_PT(752) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(759) OR ROM32_INSTR_PT(763)
     OR ROM32_INSTR_PT(774) OR ROM32_INSTR_PT(787)
     OR ROM32_INSTR_PT(790) OR ROM32_INSTR_PT(792)
     OR ROM32_INSTR_PT(795) OR ROM32_INSTR_PT(801)
     OR ROM32_INSTR_PT(803) OR ROM32_INSTR_PT(805)
     OR ROM32_INSTR_PT(807) OR ROM32_INSTR_PT(812)
     OR ROM32_INSTR_PT(817) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(823) OR ROM32_INSTR_PT(829)
     OR ROM32_INSTR_PT(831) OR ROM32_INSTR_PT(845)
     OR ROM32_INSTR_PT(847) OR ROM32_INSTR_PT(851)
     OR ROM32_INSTR_PT(853) OR ROM32_INSTR_PT(854)
     OR ROM32_INSTR_PT(857) OR ROM32_INSTR_PT(869)
     OR ROM32_INSTR_PT(872) OR ROM32_INSTR_PT(878)
     OR ROM32_INSTR_PT(881));
MQQ1860:TEMPLATE(5) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(7)
     OR ROM32_INSTR_PT(9) OR ROM32_INSTR_PT(10)
     OR ROM32_INSTR_PT(12) OR ROM32_INSTR_PT(13)
     OR ROM32_INSTR_PT(14) OR ROM32_INSTR_PT(20)
     OR ROM32_INSTR_PT(26) OR ROM32_INSTR_PT(33)
     OR ROM32_INSTR_PT(37) OR ROM32_INSTR_PT(39)
     OR ROM32_INSTR_PT(41) OR ROM32_INSTR_PT(42)
     OR ROM32_INSTR_PT(45) OR ROM32_INSTR_PT(49)
     OR ROM32_INSTR_PT(51) OR ROM32_INSTR_PT(52)
     OR ROM32_INSTR_PT(53) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(59)
     OR ROM32_INSTR_PT(63) OR ROM32_INSTR_PT(66)
     OR ROM32_INSTR_PT(67) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(73) OR ROM32_INSTR_PT(83)
     OR ROM32_INSTR_PT(84) OR ROM32_INSTR_PT(85)
     OR ROM32_INSTR_PT(87) OR ROM32_INSTR_PT(90)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(96)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(102) OR ROM32_INSTR_PT(103)
     OR ROM32_INSTR_PT(106) OR ROM32_INSTR_PT(109)
     OR ROM32_INSTR_PT(110) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(124) OR ROM32_INSTR_PT(130)
     OR ROM32_INSTR_PT(131) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(139) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(142) OR ROM32_INSTR_PT(143)
     OR ROM32_INSTR_PT(144) OR ROM32_INSTR_PT(153)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(159) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(164) OR ROM32_INSTR_PT(169)
     OR ROM32_INSTR_PT(170) OR ROM32_INSTR_PT(176)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(180)
     OR ROM32_INSTR_PT(181) OR ROM32_INSTR_PT(183)
     OR ROM32_INSTR_PT(184) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(192) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(196) OR ROM32_INSTR_PT(199)
     OR ROM32_INSTR_PT(202) OR ROM32_INSTR_PT(203)
     OR ROM32_INSTR_PT(204) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(206) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(212) OR ROM32_INSTR_PT(216)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(232)
     OR ROM32_INSTR_PT(233) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(241)
     OR ROM32_INSTR_PT(243) OR ROM32_INSTR_PT(244)
     OR ROM32_INSTR_PT(249) OR ROM32_INSTR_PT(252)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(259) OR ROM32_INSTR_PT(260)
     OR ROM32_INSTR_PT(261) OR ROM32_INSTR_PT(264)
     OR ROM32_INSTR_PT(266) OR ROM32_INSTR_PT(267)
     OR ROM32_INSTR_PT(268) OR ROM32_INSTR_PT(269)
     OR ROM32_INSTR_PT(271) OR ROM32_INSTR_PT(274)
     OR ROM32_INSTR_PT(276) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(280) OR ROM32_INSTR_PT(282)
     OR ROM32_INSTR_PT(284) OR ROM32_INSTR_PT(288)
     OR ROM32_INSTR_PT(290) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(306) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(310) OR ROM32_INSTR_PT(318)
     OR ROM32_INSTR_PT(323) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(346)
     OR ROM32_INSTR_PT(348) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(353) OR ROM32_INSTR_PT(356)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(363)
     OR ROM32_INSTR_PT(364) OR ROM32_INSTR_PT(367)
     OR ROM32_INSTR_PT(371) OR ROM32_INSTR_PT(373)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(382) OR ROM32_INSTR_PT(383)
     OR ROM32_INSTR_PT(386) OR ROM32_INSTR_PT(390)
     OR ROM32_INSTR_PT(392) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(396) OR ROM32_INSTR_PT(400)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(405)
     OR ROM32_INSTR_PT(406) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(413) OR ROM32_INSTR_PT(415)
     OR ROM32_INSTR_PT(417) OR ROM32_INSTR_PT(422)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(425) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(428) OR ROM32_INSTR_PT(430)
     OR ROM32_INSTR_PT(431) OR ROM32_INSTR_PT(434)
     OR ROM32_INSTR_PT(435) OR ROM32_INSTR_PT(436)
     OR ROM32_INSTR_PT(438) OR ROM32_INSTR_PT(441)
     OR ROM32_INSTR_PT(442) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(445) OR ROM32_INSTR_PT(449)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(452)
     OR ROM32_INSTR_PT(453) OR ROM32_INSTR_PT(458)
     OR ROM32_INSTR_PT(464) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(474)
     OR ROM32_INSTR_PT(475) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(481)
     OR ROM32_INSTR_PT(482) OR ROM32_INSTR_PT(484)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(491) OR ROM32_INSTR_PT(494)
     OR ROM32_INSTR_PT(495) OR ROM32_INSTR_PT(501)
     OR ROM32_INSTR_PT(503) OR ROM32_INSTR_PT(507)
     OR ROM32_INSTR_PT(509) OR ROM32_INSTR_PT(511)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(517)
     OR ROM32_INSTR_PT(520) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(524)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(531)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(541) OR ROM32_INSTR_PT(544)
     OR ROM32_INSTR_PT(550) OR ROM32_INSTR_PT(551)
     OR ROM32_INSTR_PT(552) OR ROM32_INSTR_PT(554)
     OR ROM32_INSTR_PT(555) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(569)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(575)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(580)
     OR ROM32_INSTR_PT(581) OR ROM32_INSTR_PT(582)
     OR ROM32_INSTR_PT(583) OR ROM32_INSTR_PT(584)
     OR ROM32_INSTR_PT(588) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(601)
     OR ROM32_INSTR_PT(602) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(609) OR ROM32_INSTR_PT(610)
     OR ROM32_INSTR_PT(613) OR ROM32_INSTR_PT(615)
     OR ROM32_INSTR_PT(616) OR ROM32_INSTR_PT(617)
     OR ROM32_INSTR_PT(620) OR ROM32_INSTR_PT(622)
     OR ROM32_INSTR_PT(624) OR ROM32_INSTR_PT(626)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(634)
     OR ROM32_INSTR_PT(638) OR ROM32_INSTR_PT(639)
     OR ROM32_INSTR_PT(642) OR ROM32_INSTR_PT(643)
     OR ROM32_INSTR_PT(654) OR ROM32_INSTR_PT(660)
     OR ROM32_INSTR_PT(663) OR ROM32_INSTR_PT(664)
     OR ROM32_INSTR_PT(666) OR ROM32_INSTR_PT(674)
     OR ROM32_INSTR_PT(677) OR ROM32_INSTR_PT(684)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(693)
     OR ROM32_INSTR_PT(697) OR ROM32_INSTR_PT(708)
     OR ROM32_INSTR_PT(711) OR ROM32_INSTR_PT(713)
     OR ROM32_INSTR_PT(718) OR ROM32_INSTR_PT(719)
     OR ROM32_INSTR_PT(726) OR ROM32_INSTR_PT(729)
     OR ROM32_INSTR_PT(745) OR ROM32_INSTR_PT(755)
     OR ROM32_INSTR_PT(762) OR ROM32_INSTR_PT(763)
     OR ROM32_INSTR_PT(792) OR ROM32_INSTR_PT(805)
     OR ROM32_INSTR_PT(812) OR ROM32_INSTR_PT(818)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(829)
     OR ROM32_INSTR_PT(831) OR ROM32_INSTR_PT(845)
     OR ROM32_INSTR_PT(853) OR ROM32_INSTR_PT(854)
     OR ROM32_INSTR_PT(855) OR ROM32_INSTR_PT(857)
     OR ROM32_INSTR_PT(862) OR ROM32_INSTR_PT(870)
     OR ROM32_INSTR_PT(872) OR ROM32_INSTR_PT(878)
    );
MQQ1861:TEMPLATE(6) <= 
    ('0');
MQQ1862:TEMPLATE(7) <= 
    ('0');
MQQ1863:TEMPLATE(8) <= 
    ('0');
MQQ1864:TEMPLATE(9) <= 
    (ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(8)
     OR ROM32_INSTR_PT(10) OR ROM32_INSTR_PT(12)
     OR ROM32_INSTR_PT(14) OR ROM32_INSTR_PT(17)
     OR ROM32_INSTR_PT(23) OR ROM32_INSTR_PT(28)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(37)
     OR ROM32_INSTR_PT(42) OR ROM32_INSTR_PT(45)
     OR ROM32_INSTR_PT(53) OR ROM32_INSTR_PT(55)
     OR ROM32_INSTR_PT(56) OR ROM32_INSTR_PT(60)
     OR ROM32_INSTR_PT(63) OR ROM32_INSTR_PT(73)
     OR ROM32_INSTR_PT(74) OR ROM32_INSTR_PT(85)
     OR ROM32_INSTR_PT(87) OR ROM32_INSTR_PT(90)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(102)
     OR ROM32_INSTR_PT(103) OR ROM32_INSTR_PT(105)
     OR ROM32_INSTR_PT(106) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(120) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(130) OR ROM32_INSTR_PT(134)
     OR ROM32_INSTR_PT(135) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(142) OR ROM32_INSTR_PT(148)
     OR ROM32_INSTR_PT(154) OR ROM32_INSTR_PT(155)
     OR ROM32_INSTR_PT(162) OR ROM32_INSTR_PT(172)
     OR ROM32_INSTR_PT(174) OR ROM32_INSTR_PT(175)
     OR ROM32_INSTR_PT(176) OR ROM32_INSTR_PT(177)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(180)
     OR ROM32_INSTR_PT(181) OR ROM32_INSTR_PT(184)
     OR ROM32_INSTR_PT(187) OR ROM32_INSTR_PT(192)
     OR ROM32_INSTR_PT(193) OR ROM32_INSTR_PT(199)
     OR ROM32_INSTR_PT(202) OR ROM32_INSTR_PT(209)
     OR ROM32_INSTR_PT(214) OR ROM32_INSTR_PT(216)
     OR ROM32_INSTR_PT(218) OR ROM32_INSTR_PT(222)
     OR ROM32_INSTR_PT(223) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(232)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(240)
     OR ROM32_INSTR_PT(242) OR ROM32_INSTR_PT(244)
     OR ROM32_INSTR_PT(249) OR ROM32_INSTR_PT(255)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(258)
     OR ROM32_INSTR_PT(260) OR ROM32_INSTR_PT(269)
     OR ROM32_INSTR_PT(272) OR ROM32_INSTR_PT(273)
     OR ROM32_INSTR_PT(274) OR ROM32_INSTR_PT(275)
     OR ROM32_INSTR_PT(280) OR ROM32_INSTR_PT(282)
     OR ROM32_INSTR_PT(283) OR ROM32_INSTR_PT(287)
     OR ROM32_INSTR_PT(288) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(297)
     OR ROM32_INSTR_PT(299) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(309) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(319)
     OR ROM32_INSTR_PT(321) OR ROM32_INSTR_PT(338)
     OR ROM32_INSTR_PT(345) OR ROM32_INSTR_PT(348)
     OR ROM32_INSTR_PT(353) OR ROM32_INSTR_PT(357)
     OR ROM32_INSTR_PT(359) OR ROM32_INSTR_PT(362)
     OR ROM32_INSTR_PT(363) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(374)
     OR ROM32_INSTR_PT(377) OR ROM32_INSTR_PT(378)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(382)
     OR ROM32_INSTR_PT(383) OR ROM32_INSTR_PT(386)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(388)
     OR ROM32_INSTR_PT(391) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(395) OR ROM32_INSTR_PT(399)
     OR ROM32_INSTR_PT(400) OR ROM32_INSTR_PT(401)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(406)
     OR ROM32_INSTR_PT(409) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(416)
     OR ROM32_INSTR_PT(422) OR ROM32_INSTR_PT(423)
     OR ROM32_INSTR_PT(431) OR ROM32_INSTR_PT(433)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(436)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(464) OR ROM32_INSTR_PT(467)
     OR ROM32_INSTR_PT(469) OR ROM32_INSTR_PT(471)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(475)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(482)
     OR ROM32_INSTR_PT(489) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(491) OR ROM32_INSTR_PT(494)
     OR ROM32_INSTR_PT(497) OR ROM32_INSTR_PT(498)
     OR ROM32_INSTR_PT(501) OR ROM32_INSTR_PT(502)
     OR ROM32_INSTR_PT(504) OR ROM32_INSTR_PT(506)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(516)
     OR ROM32_INSTR_PT(517) OR ROM32_INSTR_PT(519)
     OR ROM32_INSTR_PT(520) OR ROM32_INSTR_PT(532)
     OR ROM32_INSTR_PT(534) OR ROM32_INSTR_PT(535)
     OR ROM32_INSTR_PT(543) OR ROM32_INSTR_PT(544)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(550)
     OR ROM32_INSTR_PT(552) OR ROM32_INSTR_PT(556)
     OR ROM32_INSTR_PT(557) OR ROM32_INSTR_PT(568)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(571)
     OR ROM32_INSTR_PT(574) OR ROM32_INSTR_PT(575)
     OR ROM32_INSTR_PT(586) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(589) OR ROM32_INSTR_PT(590)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(602)
     OR ROM32_INSTR_PT(604) OR ROM32_INSTR_PT(606)
     OR ROM32_INSTR_PT(609) OR ROM32_INSTR_PT(611)
     OR ROM32_INSTR_PT(612) OR ROM32_INSTR_PT(613)
     OR ROM32_INSTR_PT(621) OR ROM32_INSTR_PT(625)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(639)
     OR ROM32_INSTR_PT(640) OR ROM32_INSTR_PT(646)
     OR ROM32_INSTR_PT(647) OR ROM32_INSTR_PT(652)
     OR ROM32_INSTR_PT(659) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(666) OR ROM32_INSTR_PT(677)
     OR ROM32_INSTR_PT(689) OR ROM32_INSTR_PT(690)
     OR ROM32_INSTR_PT(698) OR ROM32_INSTR_PT(700)
     OR ROM32_INSTR_PT(733) OR ROM32_INSTR_PT(745)
     OR ROM32_INSTR_PT(751) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(790) OR ROM32_INSTR_PT(807)
     OR ROM32_INSTR_PT(823) OR ROM32_INSTR_PT(845)
    );
MQQ1865:TEMPLATE(10) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(13)
     OR ROM32_INSTR_PT(14) OR ROM32_INSTR_PT(16)
     OR ROM32_INSTR_PT(18) OR ROM32_INSTR_PT(32)
     OR ROM32_INSTR_PT(38) OR ROM32_INSTR_PT(41)
     OR ROM32_INSTR_PT(42) OR ROM32_INSTR_PT(45)
     OR ROM32_INSTR_PT(51) OR ROM32_INSTR_PT(52)
     OR ROM32_INSTR_PT(53) OR ROM32_INSTR_PT(57)
     OR ROM32_INSTR_PT(76) OR ROM32_INSTR_PT(77)
     OR ROM32_INSTR_PT(85) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(99) OR ROM32_INSTR_PT(113)
     OR ROM32_INSTR_PT(114) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(123)
     OR ROM32_INSTR_PT(125) OR ROM32_INSTR_PT(127)
     OR ROM32_INSTR_PT(128) OR ROM32_INSTR_PT(130)
     OR ROM32_INSTR_PT(138) OR ROM32_INSTR_PT(139)
     OR ROM32_INSTR_PT(142) OR ROM32_INSTR_PT(143)
     OR ROM32_INSTR_PT(153) OR ROM32_INSTR_PT(169)
     OR ROM32_INSTR_PT(171) OR ROM32_INSTR_PT(173)
     OR ROM32_INSTR_PT(174) OR ROM32_INSTR_PT(180)
     OR ROM32_INSTR_PT(181) OR ROM32_INSTR_PT(183)
     OR ROM32_INSTR_PT(189) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(200) OR ROM32_INSTR_PT(203)
     OR ROM32_INSTR_PT(204) OR ROM32_INSTR_PT(214)
     OR ROM32_INSTR_PT(219) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(235) OR ROM32_INSTR_PT(237)
     OR ROM32_INSTR_PT(240) OR ROM32_INSTR_PT(241)
     OR ROM32_INSTR_PT(250) OR ROM32_INSTR_PT(251)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(261) OR ROM32_INSTR_PT(267)
     OR ROM32_INSTR_PT(270) OR ROM32_INSTR_PT(271)
     OR ROM32_INSTR_PT(274) OR ROM32_INSTR_PT(276)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(328) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(363)
     OR ROM32_INSTR_PT(364) OR ROM32_INSTR_PT(365)
     OR ROM32_INSTR_PT(370) OR ROM32_INSTR_PT(371)
     OR ROM32_INSTR_PT(376) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(390) OR ROM32_INSTR_PT(395)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(400)
     OR ROM32_INSTR_PT(404) OR ROM32_INSTR_PT(418)
     OR ROM32_INSTR_PT(419) OR ROM32_INSTR_PT(421)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(439)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(446)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(468)
     OR ROM32_INSTR_PT(473) OR ROM32_INSTR_PT(477)
     OR ROM32_INSTR_PT(478) OR ROM32_INSTR_PT(480)
     OR ROM32_INSTR_PT(489) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(504) OR ROM32_INSTR_PT(505)
     OR ROM32_INSTR_PT(508) OR ROM32_INSTR_PT(509)
     OR ROM32_INSTR_PT(517) OR ROM32_INSTR_PT(524)
     OR ROM32_INSTR_PT(527) OR ROM32_INSTR_PT(531)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(537)
     OR ROM32_INSTR_PT(538) OR ROM32_INSTR_PT(546)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(555)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(562)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(578)
     OR ROM32_INSTR_PT(582) OR ROM32_INSTR_PT(585)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(593)
     OR ROM32_INSTR_PT(595) OR ROM32_INSTR_PT(597)
     OR ROM32_INSTR_PT(598) OR ROM32_INSTR_PT(603)
     OR ROM32_INSTR_PT(608) OR ROM32_INSTR_PT(615)
     OR ROM32_INSTR_PT(624) OR ROM32_INSTR_PT(626)
     OR ROM32_INSTR_PT(629) OR ROM32_INSTR_PT(635)
     OR ROM32_INSTR_PT(641) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(654)
     OR ROM32_INSTR_PT(680) OR ROM32_INSTR_PT(683)
     OR ROM32_INSTR_PT(689) OR ROM32_INSTR_PT(708)
     OR ROM32_INSTR_PT(713) OR ROM32_INSTR_PT(718)
     OR ROM32_INSTR_PT(720) OR ROM32_INSTR_PT(728)
     OR ROM32_INSTR_PT(729) OR ROM32_INSTR_PT(731)
     OR ROM32_INSTR_PT(755) OR ROM32_INSTR_PT(763)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(857)
     OR ROM32_INSTR_PT(872));
MQQ1866:TEMPLATE(11) <= 
    ('0');
MQQ1867:TEMPLATE(12) <= 
    ('0');
MQQ1868:TEMPLATE(13) <= 
    ('0');
MQQ1869:TEMPLATE(14) <= 
    (ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(10)
     OR ROM32_INSTR_PT(12) OR ROM32_INSTR_PT(14)
     OR ROM32_INSTR_PT(16) OR ROM32_INSTR_PT(20)
     OR ROM32_INSTR_PT(23) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(32) OR ROM32_INSTR_PT(34)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(37)
     OR ROM32_INSTR_PT(42) OR ROM32_INSTR_PT(52)
     OR ROM32_INSTR_PT(53) OR ROM32_INSTR_PT(55)
     OR ROM32_INSTR_PT(56) OR ROM32_INSTR_PT(63)
     OR ROM32_INSTR_PT(67) OR ROM32_INSTR_PT(73)
     OR ROM32_INSTR_PT(77) OR ROM32_INSTR_PT(79)
     OR ROM32_INSTR_PT(85) OR ROM32_INSTR_PT(87)
     OR ROM32_INSTR_PT(90) OR ROM32_INSTR_PT(92)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(99) OR ROM32_INSTR_PT(103)
     OR ROM32_INSTR_PT(105) OR ROM32_INSTR_PT(111)
     OR ROM32_INSTR_PT(114) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(125) OR ROM32_INSTR_PT(127)
     OR ROM32_INSTR_PT(130) OR ROM32_INSTR_PT(138)
     OR ROM32_INSTR_PT(143) OR ROM32_INSTR_PT(155)
     OR ROM32_INSTR_PT(169) OR ROM32_INSTR_PT(171)
     OR ROM32_INSTR_PT(172) OR ROM32_INSTR_PT(174)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(181)
     OR ROM32_INSTR_PT(184) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(196) OR ROM32_INSTR_PT(200)
     OR ROM32_INSTR_PT(202) OR ROM32_INSTR_PT(209)
     OR ROM32_INSTR_PT(214) OR ROM32_INSTR_PT(216)
     OR ROM32_INSTR_PT(218) OR ROM32_INSTR_PT(219)
     OR ROM32_INSTR_PT(224) OR ROM32_INSTR_PT(227)
     OR ROM32_INSTR_PT(229) OR ROM32_INSTR_PT(232)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(240)
     OR ROM32_INSTR_PT(250) OR ROM32_INSTR_PT(257)
     OR ROM32_INSTR_PT(259) OR ROM32_INSTR_PT(261)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(267)
     OR ROM32_INSTR_PT(269) OR ROM32_INSTR_PT(270)
     OR ROM32_INSTR_PT(271) OR ROM32_INSTR_PT(272)
     OR ROM32_INSTR_PT(273) OR ROM32_INSTR_PT(274)
     OR ROM32_INSTR_PT(275) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(280) OR ROM32_INSTR_PT(283)
     OR ROM32_INSTR_PT(284) OR ROM32_INSTR_PT(288)
     OR ROM32_INSTR_PT(290) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(299) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(309) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(321) OR ROM32_INSTR_PT(328)
     OR ROM32_INSTR_PT(345) OR ROM32_INSTR_PT(348)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(362)
     OR ROM32_INSTR_PT(363) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(368)
     OR ROM32_INSTR_PT(370) OR ROM32_INSTR_PT(371)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(383)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(390)
     OR ROM32_INSTR_PT(392) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(395) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(400) OR ROM32_INSTR_PT(401)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(406)
     OR ROM32_INSTR_PT(411) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(418) OR ROM32_INSTR_PT(421)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(433) OR ROM32_INSTR_PT(436)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(445)
     OR ROM32_INSTR_PT(449) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(456) OR ROM32_INSTR_PT(464)
     OR ROM32_INSTR_PT(469) OR ROM32_INSTR_PT(472)
     OR ROM32_INSTR_PT(475) OR ROM32_INSTR_PT(476)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(480)
     OR ROM32_INSTR_PT(481) OR ROM32_INSTR_PT(482)
     OR ROM32_INSTR_PT(484) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(494) OR ROM32_INSTR_PT(497)
     OR ROM32_INSTR_PT(502) OR ROM32_INSTR_PT(508)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(517)
     OR ROM32_INSTR_PT(519) OR ROM32_INSTR_PT(520)
     OR ROM32_INSTR_PT(521) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(524) OR ROM32_INSTR_PT(532)
     OR ROM32_INSTR_PT(534) OR ROM32_INSTR_PT(535)
     OR ROM32_INSTR_PT(536) OR ROM32_INSTR_PT(541)
     OR ROM32_INSTR_PT(543) OR ROM32_INSTR_PT(546)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(550)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(556)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(565)
     OR ROM32_INSTR_PT(568) OR ROM32_INSTR_PT(570)
     OR ROM32_INSTR_PT(574) OR ROM32_INSTR_PT(575)
     OR ROM32_INSTR_PT(578) OR ROM32_INSTR_PT(582)
     OR ROM32_INSTR_PT(585) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(590) OR ROM32_INSTR_PT(595)
     OR ROM32_INSTR_PT(602) OR ROM32_INSTR_PT(603)
     OR ROM32_INSTR_PT(606) OR ROM32_INSTR_PT(607)
     OR ROM32_INSTR_PT(611) OR ROM32_INSTR_PT(612)
     OR ROM32_INSTR_PT(617) OR ROM32_INSTR_PT(621)
     OR ROM32_INSTR_PT(625) OR ROM32_INSTR_PT(630)
     OR ROM32_INSTR_PT(633) OR ROM32_INSTR_PT(635)
     OR ROM32_INSTR_PT(639) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(647)
     OR ROM32_INSTR_PT(666) OR ROM32_INSTR_PT(677)
     OR ROM32_INSTR_PT(680) OR ROM32_INSTR_PT(689)
     OR ROM32_INSTR_PT(690) OR ROM32_INSTR_PT(698)
     OR ROM32_INSTR_PT(718) OR ROM32_INSTR_PT(731)
     OR ROM32_INSTR_PT(736) OR ROM32_INSTR_PT(745)
     OR ROM32_INSTR_PT(755) OR ROM32_INSTR_PT(762)
     OR ROM32_INSTR_PT(770) OR ROM32_INSTR_PT(818)
     OR ROM32_INSTR_PT(855) OR ROM32_INSTR_PT(862)
     OR ROM32_INSTR_PT(870));
MQQ1870:TEMPLATE(15) <= 
    (ROM32_INSTR_PT(8) OR ROM32_INSTR_PT(14)
     OR ROM32_INSTR_PT(17) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(34) OR ROM32_INSTR_PT(53)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(74)
     OR ROM32_INSTR_PT(79) OR ROM32_INSTR_PT(84)
     OR ROM32_INSTR_PT(92) OR ROM32_INSTR_PT(102)
     OR ROM32_INSTR_PT(111) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(117) OR ROM32_INSTR_PT(122)
     OR ROM32_INSTR_PT(123) OR ROM32_INSTR_PT(134)
     OR ROM32_INSTR_PT(141) OR ROM32_INSTR_PT(148)
     OR ROM32_INSTR_PT(159) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(170) OR ROM32_INSTR_PT(173)
     OR ROM32_INSTR_PT(174) OR ROM32_INSTR_PT(203)
     OR ROM32_INSTR_PT(212) OR ROM32_INSTR_PT(214)
     OR ROM32_INSTR_PT(215) OR ROM32_INSTR_PT(220)
     OR ROM32_INSTR_PT(223) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(240) OR ROM32_INSTR_PT(259)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(271)
     OR ROM32_INSTR_PT(276) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(290) OR ROM32_INSTR_PT(294)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(301)
     OR ROM32_INSTR_PT(309) OR ROM32_INSTR_PT(346)
     OR ROM32_INSTR_PT(350) OR ROM32_INSTR_PT(356)
     OR ROM32_INSTR_PT(360) OR ROM32_INSTR_PT(368)
     OR ROM32_INSTR_PT(376) OR ROM32_INSTR_PT(382)
     OR ROM32_INSTR_PT(386) OR ROM32_INSTR_PT(392)
     OR ROM32_INSTR_PT(395) OR ROM32_INSTR_PT(404)
     OR ROM32_INSTR_PT(413) OR ROM32_INSTR_PT(422)
     OR ROM32_INSTR_PT(430) OR ROM32_INSTR_PT(431)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(438)
     OR ROM32_INSTR_PT(439) OR ROM32_INSTR_PT(442)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(459)
     OR ROM32_INSTR_PT(471) OR ROM32_INSTR_PT(474)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(477)
     OR ROM32_INSTR_PT(503) OR ROM32_INSTR_PT(505)
     OR ROM32_INSTR_PT(506) OR ROM32_INSTR_PT(517)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(532)
     OR ROM32_INSTR_PT(536) OR ROM32_INSTR_PT(538)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(580) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(593) OR ROM32_INSTR_PT(598)
     OR ROM32_INSTR_PT(599) OR ROM32_INSTR_PT(607)
     OR ROM32_INSTR_PT(608) OR ROM32_INSTR_PT(620)
     OR ROM32_INSTR_PT(659) OR ROM32_INSTR_PT(664)
     OR ROM32_INSTR_PT(689) OR ROM32_INSTR_PT(692)
     OR ROM32_INSTR_PT(711) OR ROM32_INSTR_PT(726)
     OR ROM32_INSTR_PT(829) OR ROM32_INSTR_PT(831)
     OR ROM32_INSTR_PT(845) OR ROM32_INSTR_PT(853)
    );
MQQ1871:TEMPLATE(16) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(9)
     OR ROM32_INSTR_PT(16) OR ROM32_INSTR_PT(18)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(32) OR ROM32_INSTR_PT(34)
     OR ROM32_INSTR_PT(38) OR ROM32_INSTR_PT(49)
     OR ROM32_INSTR_PT(55) OR ROM32_INSTR_PT(67)
     OR ROM32_INSTR_PT(77) OR ROM32_INSTR_PT(79)
     OR ROM32_INSTR_PT(84) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(99) OR ROM32_INSTR_PT(105)
     OR ROM32_INSTR_PT(111) OR ROM32_INSTR_PT(114)
     OR ROM32_INSTR_PT(115) OR ROM32_INSTR_PT(118)
     OR ROM32_INSTR_PT(119) OR ROM32_INSTR_PT(122)
     OR ROM32_INSTR_PT(127) OR ROM32_INSTR_PT(171)
     OR ROM32_INSTR_PT(186) OR ROM32_INSTR_PT(189)
     OR ROM32_INSTR_PT(200) OR ROM32_INSTR_PT(209)
     OR ROM32_INSTR_PT(215) OR ROM32_INSTR_PT(219)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(250)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(259)
     OR ROM32_INSTR_PT(261) OR ROM32_INSTR_PT(262)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(267)
     OR ROM32_INSTR_PT(272) OR ROM32_INSTR_PT(273)
     OR ROM32_INSTR_PT(278) OR ROM32_INSTR_PT(281)
     OR ROM32_INSTR_PT(283) OR ROM32_INSTR_PT(301)
     OR ROM32_INSTR_PT(313) OR ROM32_INSTR_PT(321)
     OR ROM32_INSTR_PT(328) OR ROM32_INSTR_PT(345)
     OR ROM32_INSTR_PT(360) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(368) OR ROM32_INSTR_PT(371)
     OR ROM32_INSTR_PT(390) OR ROM32_INSTR_PT(392)
     OR ROM32_INSTR_PT(396) OR ROM32_INSTR_PT(398)
     OR ROM32_INSTR_PT(401) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(424) OR ROM32_INSTR_PT(433)
     OR ROM32_INSTR_PT(446) OR ROM32_INSTR_PT(468)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(502) OR ROM32_INSTR_PT(519)
     OR ROM32_INSTR_PT(521) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(524) OR ROM32_INSTR_PT(537)
     OR ROM32_INSTR_PT(539) OR ROM32_INSTR_PT(554)
     OR ROM32_INSTR_PT(556) OR ROM32_INSTR_PT(562)
     OR ROM32_INSTR_PT(568) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(583) OR ROM32_INSTR_PT(590)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(595)
     OR ROM32_INSTR_PT(602) OR ROM32_INSTR_PT(607)
     OR ROM32_INSTR_PT(612) OR ROM32_INSTR_PT(614)
     OR ROM32_INSTR_PT(626) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(736)
     OR ROM32_INSTR_PT(762) OR ROM32_INSTR_PT(770)
     OR ROM32_INSTR_PT(870));
MQQ1872:TEMPLATE(17) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(16)
     OR ROM32_INSTR_PT(18) OR ROM32_INSTR_PT(20)
     OR ROM32_INSTR_PT(26) OR ROM32_INSTR_PT(32)
     OR ROM32_INSTR_PT(34) OR ROM32_INSTR_PT(37)
     OR ROM32_INSTR_PT(38) OR ROM32_INSTR_PT(43)
     OR ROM32_INSTR_PT(49) OR ROM32_INSTR_PT(55)
     OR ROM32_INSTR_PT(63) OR ROM32_INSTR_PT(73)
     OR ROM32_INSTR_PT(79) OR ROM32_INSTR_PT(80)
     OR ROM32_INSTR_PT(87) OR ROM32_INSTR_PT(90)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(99)
     OR ROM32_INSTR_PT(103) OR ROM32_INSTR_PT(105)
     OR ROM32_INSTR_PT(112) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(122) OR ROM32_INSTR_PT(127)
     OR ROM32_INSTR_PT(173) OR ROM32_INSTR_PT(184)
     OR ROM32_INSTR_PT(186) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(189) OR ROM32_INSTR_PT(200)
     OR ROM32_INSTR_PT(209) OR ROM32_INSTR_PT(216)
     OR ROM32_INSTR_PT(224) OR ROM32_INSTR_PT(227)
     OR ROM32_INSTR_PT(232) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(250)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(259)
     OR ROM32_INSTR_PT(262) OR ROM32_INSTR_PT(264)
     OR ROM32_INSTR_PT(269) OR ROM32_INSTR_PT(270)
     OR ROM32_INSTR_PT(272) OR ROM32_INSTR_PT(275)
     OR ROM32_INSTR_PT(278) OR ROM32_INSTR_PT(280)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(283)
     OR ROM32_INSTR_PT(284) OR ROM32_INSTR_PT(288)
     OR ROM32_INSTR_PT(299) OR ROM32_INSTR_PT(301)
     OR ROM32_INSTR_PT(303) OR ROM32_INSTR_PT(321)
     OR ROM32_INSTR_PT(326) OR ROM32_INSTR_PT(328)
     OR ROM32_INSTR_PT(340) OR ROM32_INSTR_PT(345)
     OR ROM32_INSTR_PT(348) OR ROM32_INSTR_PT(361)
     OR ROM32_INSTR_PT(366) OR ROM32_INSTR_PT(378)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(383)
     OR ROM32_INSTR_PT(392) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(404)
     OR ROM32_INSTR_PT(406) OR ROM32_INSTR_PT(416)
     OR ROM32_INSTR_PT(418) OR ROM32_INSTR_PT(419)
     OR ROM32_INSTR_PT(421) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(446) OR ROM32_INSTR_PT(468)
     OR ROM32_INSTR_PT(475) OR ROM32_INSTR_PT(476)
     OR ROM32_INSTR_PT(477) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(480)
     OR ROM32_INSTR_PT(481) OR ROM32_INSTR_PT(482)
     OR ROM32_INSTR_PT(490) OR ROM32_INSTR_PT(494)
     OR ROM32_INSTR_PT(497) OR ROM32_INSTR_PT(505)
     OR ROM32_INSTR_PT(508) OR ROM32_INSTR_PT(520)
     OR ROM32_INSTR_PT(521) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(534) OR ROM32_INSTR_PT(535)
     OR ROM32_INSTR_PT(537) OR ROM32_INSTR_PT(538)
     OR ROM32_INSTR_PT(546) OR ROM32_INSTR_PT(547)
     OR ROM32_INSTR_PT(550) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(562)
     OR ROM32_INSTR_PT(574) OR ROM32_INSTR_PT(578)
     OR ROM32_INSTR_PT(582) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(585) OR ROM32_INSTR_PT(591)
     OR ROM32_INSTR_PT(593) OR ROM32_INSTR_PT(598)
     OR ROM32_INSTR_PT(602) OR ROM32_INSTR_PT(606)
     OR ROM32_INSTR_PT(607) OR ROM32_INSTR_PT(608)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(635)
     OR ROM32_INSTR_PT(639) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(647)
     OR ROM32_INSTR_PT(666) OR ROM32_INSTR_PT(677)
     OR ROM32_INSTR_PT(680) OR ROM32_INSTR_PT(698)
     OR ROM32_INSTR_PT(870));
MQQ1873:TEMPLATE(18) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(18)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(34) OR ROM32_INSTR_PT(38)
     OR ROM32_INSTR_PT(49) OR ROM32_INSTR_PT(79)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(111) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(172) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(259)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(396) OR ROM32_INSTR_PT(398)
     OR ROM32_INSTR_PT(424) OR ROM32_INSTR_PT(468)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(537)
     OR ROM32_INSTR_PT(543) OR ROM32_INSTR_PT(554)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(720) OR ROM32_INSTR_PT(807)
     OR ROM32_INSTR_PT(823));
MQQ1874:TEMPLATE(19) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(14)
     OR ROM32_INSTR_PT(18) OR ROM32_INSTR_PT(20)
     OR ROM32_INSTR_PT(23) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(34) OR ROM32_INSTR_PT(38)
     OR ROM32_INSTR_PT(39) OR ROM32_INSTR_PT(42)
     OR ROM32_INSTR_PT(45) OR ROM32_INSTR_PT(49)
     OR ROM32_INSTR_PT(53) OR ROM32_INSTR_PT(57)
     OR ROM32_INSTR_PT(79) OR ROM32_INSTR_PT(85)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(101) OR ROM32_INSTR_PT(102)
     OR ROM32_INSTR_PT(110) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(141) OR ROM32_INSTR_PT(143)
     OR ROM32_INSTR_PT(144) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(178) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(203) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(206) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(232) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(243) OR ROM32_INSTR_PT(251)
     OR ROM32_INSTR_PT(252) OR ROM32_INSTR_PT(258)
     OR ROM32_INSTR_PT(268) OR ROM32_INSTR_PT(271)
     OR ROM32_INSTR_PT(278) OR ROM32_INSTR_PT(281)
     OR ROM32_INSTR_PT(289) OR ROM32_INSTR_PT(294)
     OR ROM32_INSTR_PT(306) OR ROM32_INSTR_PT(323)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(378) OR ROM32_INSTR_PT(382)
     OR ROM32_INSTR_PT(385) OR ROM32_INSTR_PT(386)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(405)
     OR ROM32_INSTR_PT(416) OR ROM32_INSTR_PT(417)
     OR ROM32_INSTR_PT(419) OR ROM32_INSTR_PT(422)
     OR ROM32_INSTR_PT(424) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(435) OR ROM32_INSTR_PT(436)
     OR ROM32_INSTR_PT(452) OR ROM32_INSTR_PT(458)
     OR ROM32_INSTR_PT(468) OR ROM32_INSTR_PT(476)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(507) OR ROM32_INSTR_PT(517)
     OR ROM32_INSTR_PT(521) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(532)
     OR ROM32_INSTR_PT(537) OR ROM32_INSTR_PT(541)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(554)
     OR ROM32_INSTR_PT(569) OR ROM32_INSTR_PT(579)
     OR ROM32_INSTR_PT(581) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(610) OR ROM32_INSTR_PT(615)
     OR ROM32_INSTR_PT(616) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(643) OR ROM32_INSTR_PT(674)
     OR ROM32_INSTR_PT(684) OR ROM32_INSTR_PT(720)
     OR ROM32_INSTR_PT(729) OR ROM32_INSTR_PT(763)
     OR ROM32_INSTR_PT(807) OR ROM32_INSTR_PT(812)
     OR ROM32_INSTR_PT(818) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(823) OR ROM32_INSTR_PT(878)
    );
MQQ1875:TEMPLATE(20) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(12)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(33)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(38)
     OR ROM32_INSTR_PT(42) OR ROM32_INSTR_PT(45)
     OR ROM32_INSTR_PT(49) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(102)
     OR ROM32_INSTR_PT(119) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(196) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(218) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(257)
     OR ROM32_INSTR_PT(258) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(306)
     OR ROM32_INSTR_PT(323) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(362) OR ROM32_INSTR_PT(367)
     OR ROM32_INSTR_PT(382) OR ROM32_INSTR_PT(386)
     OR ROM32_INSTR_PT(387) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(396) OR ROM32_INSTR_PT(398)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(422)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(431) OR ROM32_INSTR_PT(435)
     OR ROM32_INSTR_PT(452) OR ROM32_INSTR_PT(454)
     OR ROM32_INSTR_PT(456) OR ROM32_INSTR_PT(464)
     OR ROM32_INSTR_PT(469) OR ROM32_INSTR_PT(472)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(484)
     OR ROM32_INSTR_PT(504) OR ROM32_INSTR_PT(514)
     OR ROM32_INSTR_PT(516) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(537)
     OR ROM32_INSTR_PT(541) OR ROM32_INSTR_PT(543)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(577) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(584) OR ROM32_INSTR_PT(591)
     OR ROM32_INSTR_PT(611) OR ROM32_INSTR_PT(615)
     OR ROM32_INSTR_PT(625) OR ROM32_INSTR_PT(634)
     OR ROM32_INSTR_PT(638) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(684) OR ROM32_INSTR_PT(690)
     OR ROM32_INSTR_PT(718) OR ROM32_INSTR_PT(728)
     OR ROM32_INSTR_PT(751) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(763) OR ROM32_INSTR_PT(805)
     OR ROM32_INSTR_PT(818));
MQQ1876:TEMPLATE(21) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(8) OR ROM32_INSTR_PT(9)
     OR ROM32_INSTR_PT(10) OR ROM32_INSTR_PT(17)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(23)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(38)
     OR ROM32_INSTR_PT(43) OR ROM32_INSTR_PT(60)
     OR ROM32_INSTR_PT(73) OR ROM32_INSTR_PT(74)
     OR ROM32_INSTR_PT(78) OR ROM32_INSTR_PT(80)
     OR ROM32_INSTR_PT(84) OR ROM32_INSTR_PT(87)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(97) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(134) OR ROM32_INSTR_PT(148)
     OR ROM32_INSTR_PT(154) OR ROM32_INSTR_PT(172)
     OR ROM32_INSTR_PT(178) OR ROM32_INSTR_PT(179)
     OR ROM32_INSTR_PT(186) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(194) OR ROM32_INSTR_PT(202)
     OR ROM32_INSTR_PT(206) OR ROM32_INSTR_PT(215)
     OR ROM32_INSTR_PT(218) OR ROM32_INSTR_PT(223)
     OR ROM32_INSTR_PT(224) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(232) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(244) OR ROM32_INSTR_PT(251)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(261)
     OR ROM32_INSTR_PT(262) OR ROM32_INSTR_PT(267)
     OR ROM32_INSTR_PT(270) OR ROM32_INSTR_PT(273)
     OR ROM32_INSTR_PT(275) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(295) OR ROM32_INSTR_PT(297)
     OR ROM32_INSTR_PT(310) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(360)
     OR ROM32_INSTR_PT(362) OR ROM32_INSTR_PT(368)
     OR ROM32_INSTR_PT(371) OR ROM32_INSTR_PT(378)
     OR ROM32_INSTR_PT(385) OR ROM32_INSTR_PT(387)
     OR ROM32_INSTR_PT(390) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(401)
     OR ROM32_INSTR_PT(411) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(416) OR ROM32_INSTR_PT(419)
     OR ROM32_INSTR_PT(421) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(426) OR ROM32_INSTR_PT(433)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(496) OR ROM32_INSTR_PT(502)
     OR ROM32_INSTR_PT(506) OR ROM32_INSTR_PT(507)
     OR ROM32_INSTR_PT(508) OR ROM32_INSTR_PT(516)
     OR ROM32_INSTR_PT(519) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(524) OR ROM32_INSTR_PT(530)
     OR ROM32_INSTR_PT(531) OR ROM32_INSTR_PT(535)
     OR ROM32_INSTR_PT(537) OR ROM32_INSTR_PT(539)
     OR ROM32_INSTR_PT(543) OR ROM32_INSTR_PT(547)
     OR ROM32_INSTR_PT(556) OR ROM32_INSTR_PT(558)
     OR ROM32_INSTR_PT(568) OR ROM32_INSTR_PT(569)
     OR ROM32_INSTR_PT(574) OR ROM32_INSTR_PT(575)
     OR ROM32_INSTR_PT(578) OR ROM32_INSTR_PT(579)
     OR ROM32_INSTR_PT(583) OR ROM32_INSTR_PT(585)
     OR ROM32_INSTR_PT(588) OR ROM32_INSTR_PT(590)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(611)
     OR ROM32_INSTR_PT(612) OR ROM32_INSTR_PT(614)
     OR ROM32_INSTR_PT(621) OR ROM32_INSTR_PT(625)
     OR ROM32_INSTR_PT(626) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(751)
     OR ROM32_INSTR_PT(753) OR ROM32_INSTR_PT(817)
    );
MQQ1877:TEMPLATE(22) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(7)
     OR ROM32_INSTR_PT(8) OR ROM32_INSTR_PT(10)
     OR ROM32_INSTR_PT(12) OR ROM32_INSTR_PT(14)
     OR ROM32_INSTR_PT(17) OR ROM32_INSTR_PT(20)
     OR ROM32_INSTR_PT(23) OR ROM32_INSTR_PT(29)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(38)
     OR ROM32_INSTR_PT(43) OR ROM32_INSTR_PT(53)
     OR ROM32_INSTR_PT(56) OR ROM32_INSTR_PT(57)
     OR ROM32_INSTR_PT(74) OR ROM32_INSTR_PT(78)
     OR ROM32_INSTR_PT(80) OR ROM32_INSTR_PT(93)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(101) OR ROM32_INSTR_PT(114)
     OR ROM32_INSTR_PT(119) OR ROM32_INSTR_PT(122)
     OR ROM32_INSTR_PT(131) OR ROM32_INSTR_PT(134)
     OR ROM32_INSTR_PT(143) OR ROM32_INSTR_PT(148)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(163) OR ROM32_INSTR_PT(164)
     OR ROM32_INSTR_PT(171) OR ROM32_INSTR_PT(172)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(186)
     OR ROM32_INSTR_PT(196) OR ROM32_INSTR_PT(202)
     OR ROM32_INSTR_PT(203) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(207) OR ROM32_INSTR_PT(212)
     OR ROM32_INSTR_PT(218) OR ROM32_INSTR_PT(220)
     OR ROM32_INSTR_PT(223) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(229) OR ROM32_INSTR_PT(243)
     OR ROM32_INSTR_PT(244) OR ROM32_INSTR_PT(251)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(262)
     OR ROM32_INSTR_PT(271) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(295) OR ROM32_INSTR_PT(297)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(310)
     OR ROM32_INSTR_PT(323) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(362) OR ROM32_INSTR_PT(367)
     OR ROM32_INSTR_PT(376) OR ROM32_INSTR_PT(387)
     OR ROM32_INSTR_PT(392) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(396) OR ROM32_INSTR_PT(398)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(411)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(435)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(438)
     OR ROM32_INSTR_PT(452) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(456)
     OR ROM32_INSTR_PT(458) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(464) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(484) OR ROM32_INSTR_PT(486)
     OR ROM32_INSTR_PT(496) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(506) OR ROM32_INSTR_PT(511)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(516)
     OR ROM32_INSTR_PT(517) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(537)
     OR ROM32_INSTR_PT(539) OR ROM32_INSTR_PT(543)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(558)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(575)
     OR ROM32_INSTR_PT(577) OR ROM32_INSTR_PT(580)
     OR ROM32_INSTR_PT(581) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(584) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(601) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(607) OR ROM32_INSTR_PT(611)
     OR ROM32_INSTR_PT(614) OR ROM32_INSTR_PT(622)
     OR ROM32_INSTR_PT(625) OR ROM32_INSTR_PT(634)
     OR ROM32_INSTR_PT(638) OR ROM32_INSTR_PT(643)
     OR ROM32_INSTR_PT(654) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(684) OR ROM32_INSTR_PT(693)
     OR ROM32_INSTR_PT(708) OR ROM32_INSTR_PT(720)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(751)
     OR ROM32_INSTR_PT(753) OR ROM32_INSTR_PT(807)
     OR ROM32_INSTR_PT(817) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(823) OR ROM32_INSTR_PT(845)
     OR ROM32_INSTR_PT(853));
MQQ1878:TEMPLATE(23) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(12) OR ROM32_INSTR_PT(23)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(38)
     OR ROM32_INSTR_PT(56) OR ROM32_INSTR_PT(57)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(111) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(135) OR ROM32_INSTR_PT(143)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(163) OR ROM32_INSTR_PT(179)
     OR ROM32_INSTR_PT(187) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(202) OR ROM32_INSTR_PT(203)
     OR ROM32_INSTR_PT(207) OR ROM32_INSTR_PT(218)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(232) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(243) OR ROM32_INSTR_PT(244)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(254)
     OR ROM32_INSTR_PT(256) OR ROM32_INSTR_PT(257)
     OR ROM32_INSTR_PT(259) OR ROM32_INSTR_PT(260)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(275)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(282)
     OR ROM32_INSTR_PT(293) OR ROM32_INSTR_PT(310)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(362) OR ROM32_INSTR_PT(367)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(378) OR ROM32_INSTR_PT(387)
     OR ROM32_INSTR_PT(394) OR ROM32_INSTR_PT(398)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(416) OR ROM32_INSTR_PT(419)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(434)
     OR ROM32_INSTR_PT(443) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(456)
     OR ROM32_INSTR_PT(458) OR ROM32_INSTR_PT(464)
     OR ROM32_INSTR_PT(469) OR ROM32_INSTR_PT(472)
     OR ROM32_INSTR_PT(484) OR ROM32_INSTR_PT(486)
     OR ROM32_INSTR_PT(501) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(516)
     OR ROM32_INSTR_PT(531) OR ROM32_INSTR_PT(535)
     OR ROM32_INSTR_PT(537) OR ROM32_INSTR_PT(544)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(551)
     OR ROM32_INSTR_PT(557) OR ROM32_INSTR_PT(558)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(577) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(588) OR ROM32_INSTR_PT(591)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(609) OR ROM32_INSTR_PT(611)
     OR ROM32_INSTR_PT(621) OR ROM32_INSTR_PT(625)
     OR ROM32_INSTR_PT(643) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(690) OR ROM32_INSTR_PT(713)
     OR ROM32_INSTR_PT(720) OR ROM32_INSTR_PT(728)
     OR ROM32_INSTR_PT(751) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(807) OR ROM32_INSTR_PT(817)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(823)
     OR ROM32_INSTR_PT(845));
MQQ1879:TEMPLATE(24) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(4)
     OR ROM32_INSTR_PT(5) OR ROM32_INSTR_PT(10)
     OR ROM32_INSTR_PT(13) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(29) OR ROM32_INSTR_PT(34)
     OR ROM32_INSTR_PT(35) OR ROM32_INSTR_PT(41)
     OR ROM32_INSTR_PT(45) OR ROM32_INSTR_PT(51)
     OR ROM32_INSTR_PT(79) OR ROM32_INSTR_PT(93)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(100)
     OR ROM32_INSTR_PT(106) OR ROM32_INSTR_PT(116)
     OR ROM32_INSTR_PT(124) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(139) OR ROM32_INSTR_PT(142)
     OR ROM32_INSTR_PT(153) OR ROM32_INSTR_PT(159)
     OR ROM32_INSTR_PT(170) OR ROM32_INSTR_PT(172)
     OR ROM32_INSTR_PT(183) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(204) OR ROM32_INSTR_PT(218)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(241) OR ROM32_INSTR_PT(251)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(258)
     OR ROM32_INSTR_PT(260) OR ROM32_INSTR_PT(275)
     OR ROM32_INSTR_PT(276) OR ROM32_INSTR_PT(281)
     OR ROM32_INSTR_PT(282) OR ROM32_INSTR_PT(290)
     OR ROM32_INSTR_PT(293) OR ROM32_INSTR_PT(306)
     OR ROM32_INSTR_PT(309) OR ROM32_INSTR_PT(318)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(362)
     OR ROM32_INSTR_PT(363) OR ROM32_INSTR_PT(374)
     OR ROM32_INSTR_PT(385) OR ROM32_INSTR_PT(393)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(425)
     OR ROM32_INSTR_PT(426) OR ROM32_INSTR_PT(428)
     OR ROM32_INSTR_PT(430) OR ROM32_INSTR_PT(434)
     OR ROM32_INSTR_PT(437) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(454)
     OR ROM32_INSTR_PT(495) OR ROM32_INSTR_PT(501)
     OR ROM32_INSTR_PT(509) OR ROM32_INSTR_PT(516)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(531)
     OR ROM32_INSTR_PT(535) OR ROM32_INSTR_PT(543)
     OR ROM32_INSTR_PT(544) OR ROM32_INSTR_PT(547)
     OR ROM32_INSTR_PT(555) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(574) OR ROM32_INSTR_PT(575)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(587) OR ROM32_INSTR_PT(591)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(609)
     OR ROM32_INSTR_PT(611) OR ROM32_INSTR_PT(615)
     OR ROM32_INSTR_PT(621) OR ROM32_INSTR_PT(624)
     OR ROM32_INSTR_PT(625) OR ROM32_INSTR_PT(646)
     OR ROM32_INSTR_PT(663) OR ROM32_INSTR_PT(690)
     OR ROM32_INSTR_PT(700) OR ROM32_INSTR_PT(729)
     OR ROM32_INSTR_PT(745) OR ROM32_INSTR_PT(763)
     OR ROM32_INSTR_PT(817) OR ROM32_INSTR_PT(845)
    );
MQQ1880:TEMPLATE(25) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(12) OR ROM32_INSTR_PT(20)
     OR ROM32_INSTR_PT(23) OR ROM32_INSTR_PT(35)
     OR ROM32_INSTR_PT(42) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(97) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(119) OR ROM32_INSTR_PT(125)
     OR ROM32_INSTR_PT(132) OR ROM32_INSTR_PT(142)
     OR ROM32_INSTR_PT(143) OR ROM32_INSTR_PT(155)
     OR ROM32_INSTR_PT(158) OR ROM32_INSTR_PT(159)
     OR ROM32_INSTR_PT(163) OR ROM32_INSTR_PT(170)
     OR ROM32_INSTR_PT(172) OR ROM32_INSTR_PT(178)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(194) OR ROM32_INSTR_PT(196)
     OR ROM32_INSTR_PT(203) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(218) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(229) OR ROM32_INSTR_PT(232)
     OR ROM32_INSTR_PT(235) OR ROM32_INSTR_PT(243)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(257) OR ROM32_INSTR_PT(275)
     OR ROM32_INSTR_PT(276) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(290)
     OR ROM32_INSTR_PT(309) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(362) OR ROM32_INSTR_PT(363)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(378) OR ROM32_INSTR_PT(385)
     OR ROM32_INSTR_PT(394) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(402)
     OR ROM32_INSTR_PT(416) OR ROM32_INSTR_PT(419)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(426) OR ROM32_INSTR_PT(430)
     OR ROM32_INSTR_PT(442) OR ROM32_INSTR_PT(454)
     OR ROM32_INSTR_PT(456) OR ROM32_INSTR_PT(458)
     OR ROM32_INSTR_PT(464) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(474)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(484)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(504) OR ROM32_INSTR_PT(514)
     OR ROM32_INSTR_PT(521) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(531)
     OR ROM32_INSTR_PT(535) OR ROM32_INSTR_PT(541)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(551)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(555)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(575) OR ROM32_INSTR_PT(577)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(611) OR ROM32_INSTR_PT(620)
     OR ROM32_INSTR_PT(629) OR ROM32_INSTR_PT(633)
     OR ROM32_INSTR_PT(642) OR ROM32_INSTR_PT(643)
     OR ROM32_INSTR_PT(654) OR ROM32_INSTR_PT(664)
     OR ROM32_INSTR_PT(690) OR ROM32_INSTR_PT(697)
     OR ROM32_INSTR_PT(708) OR ROM32_INSTR_PT(729)
     OR ROM32_INSTR_PT(731) OR ROM32_INSTR_PT(745)
     OR ROM32_INSTR_PT(792) OR ROM32_INSTR_PT(817)
     OR ROM32_INSTR_PT(818) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(829));
MQQ1881:TEMPLATE(26) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(4)
     OR ROM32_INSTR_PT(5) OR ROM32_INSTR_PT(6)
     OR ROM32_INSTR_PT(8) OR ROM32_INSTR_PT(9)
     OR ROM32_INSTR_PT(10) OR ROM32_INSTR_PT(12)
     OR ROM32_INSTR_PT(13) OR ROM32_INSTR_PT(17)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(23)
     OR ROM32_INSTR_PT(26) OR ROM32_INSTR_PT(29)
     OR ROM32_INSTR_PT(33) OR ROM32_INSTR_PT(35)
     OR ROM32_INSTR_PT(37) OR ROM32_INSTR_PT(39)
     OR ROM32_INSTR_PT(41) OR ROM32_INSTR_PT(43)
     OR ROM32_INSTR_PT(45) OR ROM32_INSTR_PT(49)
     OR ROM32_INSTR_PT(50) OR ROM32_INSTR_PT(51)
     OR ROM32_INSTR_PT(52) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(59)
     OR ROM32_INSTR_PT(60) OR ROM32_INSTR_PT(63)
     OR ROM32_INSTR_PT(66) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(73) OR ROM32_INSTR_PT(74)
     OR ROM32_INSTR_PT(78) OR ROM32_INSTR_PT(80)
     OR ROM32_INSTR_PT(83) OR ROM32_INSTR_PT(84)
     OR ROM32_INSTR_PT(85) OR ROM32_INSTR_PT(87)
     OR ROM32_INSTR_PT(90) OR ROM32_INSTR_PT(92)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(96) OR ROM32_INSTR_PT(97)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(102) OR ROM32_INSTR_PT(103)
     OR ROM32_INSTR_PT(106) OR ROM32_INSTR_PT(109)
     OR ROM32_INSTR_PT(110) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(124) OR ROM32_INSTR_PT(130)
     OR ROM32_INSTR_PT(134) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(139) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(142) OR ROM32_INSTR_PT(143)
     OR ROM32_INSTR_PT(144) OR ROM32_INSTR_PT(148)
     OR ROM32_INSTR_PT(153) OR ROM32_INSTR_PT(154)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(159) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(169) OR ROM32_INSTR_PT(172)
     OR ROM32_INSTR_PT(174) OR ROM32_INSTR_PT(176)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(180)
     OR ROM32_INSTR_PT(181) OR ROM32_INSTR_PT(183)
     OR ROM32_INSTR_PT(184) OR ROM32_INSTR_PT(186)
     OR ROM32_INSTR_PT(192) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(196) OR ROM32_INSTR_PT(199)
     OR ROM32_INSTR_PT(202) OR ROM32_INSTR_PT(203)
     OR ROM32_INSTR_PT(204) OR ROM32_INSTR_PT(206)
     OR ROM32_INSTR_PT(207) OR ROM32_INSTR_PT(216)
     OR ROM32_INSTR_PT(218) OR ROM32_INSTR_PT(220)
     OR ROM32_INSTR_PT(223) OR ROM32_INSTR_PT(224)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(233)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(241)
     OR ROM32_INSTR_PT(243) OR ROM32_INSTR_PT(244)
     OR ROM32_INSTR_PT(249) OR ROM32_INSTR_PT(251)
     OR ROM32_INSTR_PT(252) OR ROM32_INSTR_PT(254)
     OR ROM32_INSTR_PT(256) OR ROM32_INSTR_PT(257)
     OR ROM32_INSTR_PT(259) OR ROM32_INSTR_PT(260)
     OR ROM32_INSTR_PT(261) OR ROM32_INSTR_PT(262)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(266)
     OR ROM32_INSTR_PT(267) OR ROM32_INSTR_PT(268)
     OR ROM32_INSTR_PT(269) OR ROM32_INSTR_PT(270)
     OR ROM32_INSTR_PT(273) OR ROM32_INSTR_PT(274)
     OR ROM32_INSTR_PT(275) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(280) OR ROM32_INSTR_PT(281)
     OR ROM32_INSTR_PT(282) OR ROM32_INSTR_PT(284)
     OR ROM32_INSTR_PT(288) OR ROM32_INSTR_PT(289)
     OR ROM32_INSTR_PT(290) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(306) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(310) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(346)
     OR ROM32_INSTR_PT(348) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(353) OR ROM32_INSTR_PT(356)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(362)
     OR ROM32_INSTR_PT(364) OR ROM32_INSTR_PT(367)
     OR ROM32_INSTR_PT(371) OR ROM32_INSTR_PT(373)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(382) OR ROM32_INSTR_PT(383)
     OR ROM32_INSTR_PT(386) OR ROM32_INSTR_PT(387)
     OR ROM32_INSTR_PT(390) OR ROM32_INSTR_PT(392)
     OR ROM32_INSTR_PT(394) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(400)
     OR ROM32_INSTR_PT(401) OR ROM32_INSTR_PT(402)
     OR ROM32_INSTR_PT(405) OR ROM32_INSTR_PT(406)
     OR ROM32_INSTR_PT(409) OR ROM32_INSTR_PT(411)
     OR ROM32_INSTR_PT(412) OR ROM32_INSTR_PT(415)
     OR ROM32_INSTR_PT(417) OR ROM32_INSTR_PT(421)
     OR ROM32_INSTR_PT(422) OR ROM32_INSTR_PT(423)
     OR ROM32_INSTR_PT(424) OR ROM32_INSTR_PT(425)
     OR ROM32_INSTR_PT(426) OR ROM32_INSTR_PT(428)
     OR ROM32_INSTR_PT(431) OR ROM32_INSTR_PT(433)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(437)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(454) OR ROM32_INSTR_PT(458)
     OR ROM32_INSTR_PT(459) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(464) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(475)
     OR ROM32_INSTR_PT(478) OR ROM32_INSTR_PT(479)
     OR ROM32_INSTR_PT(481) OR ROM32_INSTR_PT(482)
     OR ROM32_INSTR_PT(484) OR ROM32_INSTR_PT(486)
     OR ROM32_INSTR_PT(490) OR ROM32_INSTR_PT(491)
     OR ROM32_INSTR_PT(494) OR ROM32_INSTR_PT(495)
     OR ROM32_INSTR_PT(496) OR ROM32_INSTR_PT(501)
     OR ROM32_INSTR_PT(502) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(506) OR ROM32_INSTR_PT(507)
     OR ROM32_INSTR_PT(508) OR ROM32_INSTR_PT(509)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(516)
     OR ROM32_INSTR_PT(519) OR ROM32_INSTR_PT(520)
     OR ROM32_INSTR_PT(521) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(524) OR ROM32_INSTR_PT(530)
     OR ROM32_INSTR_PT(531) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(535) OR ROM32_INSTR_PT(539)
     OR ROM32_INSTR_PT(543) OR ROM32_INSTR_PT(544)
     OR ROM32_INSTR_PT(547) OR ROM32_INSTR_PT(550)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(555)
     OR ROM32_INSTR_PT(556) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(568) OR ROM32_INSTR_PT(569)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(575) OR ROM32_INSTR_PT(578)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(582) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(585) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(590) OR ROM32_INSTR_PT(591)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(602)
     OR ROM32_INSTR_PT(603) OR ROM32_INSTR_PT(605)
     OR ROM32_INSTR_PT(609) OR ROM32_INSTR_PT(610)
     OR ROM32_INSTR_PT(611) OR ROM32_INSTR_PT(612)
     OR ROM32_INSTR_PT(613) OR ROM32_INSTR_PT(614)
     OR ROM32_INSTR_PT(615) OR ROM32_INSTR_PT(621)
     OR ROM32_INSTR_PT(624) OR ROM32_INSTR_PT(625)
     OR ROM32_INSTR_PT(626) OR ROM32_INSTR_PT(629)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(639)
     OR ROM32_INSTR_PT(640) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(643) OR ROM32_INSTR_PT(654)
     OR ROM32_INSTR_PT(660) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(664) OR ROM32_INSTR_PT(666)
     OR ROM32_INSTR_PT(674) OR ROM32_INSTR_PT(677)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(697)
     OR ROM32_INSTR_PT(708) OR ROM32_INSTR_PT(711)
     OR ROM32_INSTR_PT(713) OR ROM32_INSTR_PT(718)
     OR ROM32_INSTR_PT(719) OR ROM32_INSTR_PT(720)
     OR ROM32_INSTR_PT(729) OR ROM32_INSTR_PT(755)
     OR ROM32_INSTR_PT(763) OR ROM32_INSTR_PT(792)
     OR ROM32_INSTR_PT(805) OR ROM32_INSTR_PT(807)
     OR ROM32_INSTR_PT(812) OR ROM32_INSTR_PT(817)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(823)
     OR ROM32_INSTR_PT(829) OR ROM32_INSTR_PT(831)
     OR ROM32_INSTR_PT(845) OR ROM32_INSTR_PT(854)
     OR ROM32_INSTR_PT(855) OR ROM32_INSTR_PT(857)
     OR ROM32_INSTR_PT(862) OR ROM32_INSTR_PT(870)
     OR ROM32_INSTR_PT(872) OR ROM32_INSTR_PT(878)
    );
MQQ1882:TEMPLATE(27) <= 
    (ROM32_INSTR_PT(4) OR ROM32_INSTR_PT(5)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(7)
     OR ROM32_INSTR_PT(8) OR ROM32_INSTR_PT(9)
     OR ROM32_INSTR_PT(10) OR ROM32_INSTR_PT(12)
     OR ROM32_INSTR_PT(14) OR ROM32_INSTR_PT(17)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(33) OR ROM32_INSTR_PT(37)
     OR ROM32_INSTR_PT(39) OR ROM32_INSTR_PT(42)
     OR ROM32_INSTR_PT(45) OR ROM32_INSTR_PT(49)
     OR ROM32_INSTR_PT(52) OR ROM32_INSTR_PT(53)
     OR ROM32_INSTR_PT(56) OR ROM32_INSTR_PT(57)
     OR ROM32_INSTR_PT(59) OR ROM32_INSTR_PT(63)
     OR ROM32_INSTR_PT(66) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(74) OR ROM32_INSTR_PT(83)
     OR ROM32_INSTR_PT(84) OR ROM32_INSTR_PT(85)
     OR ROM32_INSTR_PT(90) OR ROM32_INSTR_PT(93)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(96)
     OR ROM32_INSTR_PT(101) OR ROM32_INSTR_PT(102)
     OR ROM32_INSTR_PT(103) OR ROM32_INSTR_PT(109)
     OR ROM32_INSTR_PT(110) OR ROM32_INSTR_PT(114)
     OR ROM32_INSTR_PT(115) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(130) OR ROM32_INSTR_PT(131)
     OR ROM32_INSTR_PT(134) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(142) OR ROM32_INSTR_PT(143)
     OR ROM32_INSTR_PT(144) OR ROM32_INSTR_PT(148)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(159) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(164) OR ROM32_INSTR_PT(169)
     OR ROM32_INSTR_PT(170) OR ROM32_INSTR_PT(171)
     OR ROM32_INSTR_PT(176) OR ROM32_INSTR_PT(178)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(180)
     OR ROM32_INSTR_PT(181) OR ROM32_INSTR_PT(184)
     OR ROM32_INSTR_PT(187) OR ROM32_INSTR_PT(192)
     OR ROM32_INSTR_PT(194) OR ROM32_INSTR_PT(196)
     OR ROM32_INSTR_PT(199) OR ROM32_INSTR_PT(202)
     OR ROM32_INSTR_PT(203) OR ROM32_INSTR_PT(205)
     OR ROM32_INSTR_PT(206) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(212) OR ROM32_INSTR_PT(216)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(223)
     OR ROM32_INSTR_PT(224) OR ROM32_INSTR_PT(227)
     OR ROM32_INSTR_PT(232) OR ROM32_INSTR_PT(233)
     OR ROM32_INSTR_PT(235) OR ROM32_INSTR_PT(238)
     OR ROM32_INSTR_PT(240) OR ROM32_INSTR_PT(243)
     OR ROM32_INSTR_PT(244) OR ROM32_INSTR_PT(249)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(252)
     OR ROM32_INSTR_PT(254) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(259) OR ROM32_INSTR_PT(261)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(266)
     OR ROM32_INSTR_PT(267) OR ROM32_INSTR_PT(268)
     OR ROM32_INSTR_PT(269) OR ROM32_INSTR_PT(271)
     OR ROM32_INSTR_PT(274) OR ROM32_INSTR_PT(276)
     OR ROM32_INSTR_PT(278) OR ROM32_INSTR_PT(280)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(284)
     OR ROM32_INSTR_PT(288) OR ROM32_INSTR_PT(290)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(310) OR ROM32_INSTR_PT(323)
     OR ROM32_INSTR_PT(335) OR ROM32_INSTR_PT(344)
     OR ROM32_INSTR_PT(348) OR ROM32_INSTR_PT(350)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(363)
     OR ROM32_INSTR_PT(364) OR ROM32_INSTR_PT(367)
     OR ROM32_INSTR_PT(371) OR ROM32_INSTR_PT(373)
     OR ROM32_INSTR_PT(376) OR ROM32_INSTR_PT(378)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(382) OR ROM32_INSTR_PT(383)
     OR ROM32_INSTR_PT(386) OR ROM32_INSTR_PT(390)
     OR ROM32_INSTR_PT(392) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(395) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(400)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(405)
     OR ROM32_INSTR_PT(406) OR ROM32_INSTR_PT(411)
     OR ROM32_INSTR_PT(416) OR ROM32_INSTR_PT(417)
     OR ROM32_INSTR_PT(419) OR ROM32_INSTR_PT(422)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(424)
     OR ROM32_INSTR_PT(425) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(430) OR ROM32_INSTR_PT(431)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(435)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(438)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(442)
     OR ROM32_INSTR_PT(452) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(456) OR ROM32_INSTR_PT(458)
     OR ROM32_INSTR_PT(464) OR ROM32_INSTR_PT(469)
     OR ROM32_INSTR_PT(472) OR ROM32_INSTR_PT(474)
     OR ROM32_INSTR_PT(475) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(481)
     OR ROM32_INSTR_PT(482) OR ROM32_INSTR_PT(484)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(494)
     OR ROM32_INSTR_PT(503) OR ROM32_INSTR_PT(506)
     OR ROM32_INSTR_PT(507) OR ROM32_INSTR_PT(511)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(517)
     OR ROM32_INSTR_PT(520) OR ROM32_INSTR_PT(521)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(524)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(531)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(541) OR ROM32_INSTR_PT(550)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(555)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(569)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(575)
     OR ROM32_INSTR_PT(577) OR ROM32_INSTR_PT(579)
     OR ROM32_INSTR_PT(580) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(582) OR ROM32_INSTR_PT(583)
     OR ROM32_INSTR_PT(584) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(601) OR ROM32_INSTR_PT(602)
     OR ROM32_INSTR_PT(605) OR ROM32_INSTR_PT(610)
     OR ROM32_INSTR_PT(615) OR ROM32_INSTR_PT(620)
     OR ROM32_INSTR_PT(622) OR ROM32_INSTR_PT(626)
     OR ROM32_INSTR_PT(629) OR ROM32_INSTR_PT(630)
     OR ROM32_INSTR_PT(634) OR ROM32_INSTR_PT(638)
     OR ROM32_INSTR_PT(639) OR ROM32_INSTR_PT(640)
     OR ROM32_INSTR_PT(642) OR ROM32_INSTR_PT(643)
     OR ROM32_INSTR_PT(654) OR ROM32_INSTR_PT(660)
     OR ROM32_INSTR_PT(663) OR ROM32_INSTR_PT(664)
     OR ROM32_INSTR_PT(666) OR ROM32_INSTR_PT(674)
     OR ROM32_INSTR_PT(677) OR ROM32_INSTR_PT(684)
     OR ROM32_INSTR_PT(693) OR ROM32_INSTR_PT(697)
     OR ROM32_INSTR_PT(708) OR ROM32_INSTR_PT(719)
     OR ROM32_INSTR_PT(720) OR ROM32_INSTR_PT(729)
     OR ROM32_INSTR_PT(745) OR ROM32_INSTR_PT(755)
     OR ROM32_INSTR_PT(763) OR ROM32_INSTR_PT(792)
     OR ROM32_INSTR_PT(805) OR ROM32_INSTR_PT(807)
     OR ROM32_INSTR_PT(812) OR ROM32_INSTR_PT(818)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(823)
     OR ROM32_INSTR_PT(829) OR ROM32_INSTR_PT(831)
     OR ROM32_INSTR_PT(853) OR ROM32_INSTR_PT(854)
     OR ROM32_INSTR_PT(855) OR ROM32_INSTR_PT(862)
     OR ROM32_INSTR_PT(870) OR ROM32_INSTR_PT(878)
    );
MQQ1883:TEMPLATE(28) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(4)
     OR ROM32_INSTR_PT(5) OR ROM32_INSTR_PT(8)
     OR ROM32_INSTR_PT(9) OR ROM32_INSTR_PT(12)
     OR ROM32_INSTR_PT(13) OR ROM32_INSTR_PT(16)
     OR ROM32_INSTR_PT(17) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(32) OR ROM32_INSTR_PT(37)
     OR ROM32_INSTR_PT(39) OR ROM32_INSTR_PT(41)
     OR ROM32_INSTR_PT(45) OR ROM32_INSTR_PT(51)
     OR ROM32_INSTR_PT(52) OR ROM32_INSTR_PT(56)
     OR ROM32_INSTR_PT(57) OR ROM32_INSTR_PT(59)
     OR ROM32_INSTR_PT(63) OR ROM32_INSTR_PT(66)
     OR ROM32_INSTR_PT(67) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(73) OR ROM32_INSTR_PT(74)
     OR ROM32_INSTR_PT(77) OR ROM32_INSTR_PT(83)
     OR ROM32_INSTR_PT(84) OR ROM32_INSTR_PT(85)
     OR ROM32_INSTR_PT(87) OR ROM32_INSTR_PT(90)
     OR ROM32_INSTR_PT(93) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(98) OR ROM32_INSTR_PT(99)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(101)
     OR ROM32_INSTR_PT(102) OR ROM32_INSTR_PT(103)
     OR ROM32_INSTR_PT(106) OR ROM32_INSTR_PT(109)
     OR ROM32_INSTR_PT(114) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(118)
     OR ROM32_INSTR_PT(124) OR ROM32_INSTR_PT(125)
     OR ROM32_INSTR_PT(127) OR ROM32_INSTR_PT(132)
     OR ROM32_INSTR_PT(134) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(139) OR ROM32_INSTR_PT(141)
     OR ROM32_INSTR_PT(142) OR ROM32_INSTR_PT(143)
     OR ROM32_INSTR_PT(148) OR ROM32_INSTR_PT(153)
     OR ROM32_INSTR_PT(155) OR ROM32_INSTR_PT(158)
     OR ROM32_INSTR_PT(159) OR ROM32_INSTR_PT(163)
     OR ROM32_INSTR_PT(169) OR ROM32_INSTR_PT(171)
     OR ROM32_INSTR_PT(179) OR ROM32_INSTR_PT(183)
     OR ROM32_INSTR_PT(184) OR ROM32_INSTR_PT(192)
     OR ROM32_INSTR_PT(194) OR ROM32_INSTR_PT(196)
     OR ROM32_INSTR_PT(199) OR ROM32_INSTR_PT(200)
     OR ROM32_INSTR_PT(202) OR ROM32_INSTR_PT(203)
     OR ROM32_INSTR_PT(204) OR ROM32_INSTR_PT(207)
     OR ROM32_INSTR_PT(216) OR ROM32_INSTR_PT(219)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(223)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(238)
     OR ROM32_INSTR_PT(241) OR ROM32_INSTR_PT(243)
     OR ROM32_INSTR_PT(249) OR ROM32_INSTR_PT(250)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(254)
     OR ROM32_INSTR_PT(256) OR ROM32_INSTR_PT(259)
     OR ROM32_INSTR_PT(260) OR ROM32_INSTR_PT(261)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(266)
     OR ROM32_INSTR_PT(267) OR ROM32_INSTR_PT(268)
     OR ROM32_INSTR_PT(269) OR ROM32_INSTR_PT(270)
     OR ROM32_INSTR_PT(273) OR ROM32_INSTR_PT(280)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(282)
     OR ROM32_INSTR_PT(284) OR ROM32_INSTR_PT(288)
     OR ROM32_INSTR_PT(290) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(294) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(306) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(313) OR ROM32_INSTR_PT(318)
     OR ROM32_INSTR_PT(328) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(348)
     OR ROM32_INSTR_PT(350) OR ROM32_INSTR_PT(361)
     OR ROM32_INSTR_PT(367) OR ROM32_INSTR_PT(371)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(376)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(382) OR ROM32_INSTR_PT(383)
     OR ROM32_INSTR_PT(386) OR ROM32_INSTR_PT(390)
     OR ROM32_INSTR_PT(392) OR ROM32_INSTR_PT(394)
     OR ROM32_INSTR_PT(398) OR ROM32_INSTR_PT(401)
     OR ROM32_INSTR_PT(402) OR ROM32_INSTR_PT(406)
     OR ROM32_INSTR_PT(409) OR ROM32_INSTR_PT(411)
     OR ROM32_INSTR_PT(412) OR ROM32_INSTR_PT(415)
     OR ROM32_INSTR_PT(421) OR ROM32_INSTR_PT(422)
     OR ROM32_INSTR_PT(423) OR ROM32_INSTR_PT(425)
     OR ROM32_INSTR_PT(426) OR ROM32_INSTR_PT(428)
     OR ROM32_INSTR_PT(431) OR ROM32_INSTR_PT(433)
     OR ROM32_INSTR_PT(437) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(453)
     OR ROM32_INSTR_PT(458) OR ROM32_INSTR_PT(464)
     OR ROM32_INSTR_PT(469) OR ROM32_INSTR_PT(472)
     OR ROM32_INSTR_PT(475) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(481)
     OR ROM32_INSTR_PT(482) OR ROM32_INSTR_PT(484)
     OR ROM32_INSTR_PT(486) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(491) OR ROM32_INSTR_PT(494)
     OR ROM32_INSTR_PT(495) OR ROM32_INSTR_PT(501)
     OR ROM32_INSTR_PT(502) OR ROM32_INSTR_PT(503)
     OR ROM32_INSTR_PT(504) OR ROM32_INSTR_PT(506)
     OR ROM32_INSTR_PT(508) OR ROM32_INSTR_PT(509)
     OR ROM32_INSTR_PT(514) OR ROM32_INSTR_PT(519)
     OR ROM32_INSTR_PT(520) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(524) OR ROM32_INSTR_PT(530)
     OR ROM32_INSTR_PT(531) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(544) OR ROM32_INSTR_PT(550)
     OR ROM32_INSTR_PT(551) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(555)
     OR ROM32_INSTR_PT(556) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(568) OR ROM32_INSTR_PT(578)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(581)
     OR ROM32_INSTR_PT(582) OR ROM32_INSTR_PT(585)
     OR ROM32_INSTR_PT(588) OR ROM32_INSTR_PT(590)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(595)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(602)
     OR ROM32_INSTR_PT(605) OR ROM32_INSTR_PT(609)
     OR ROM32_INSTR_PT(612) OR ROM32_INSTR_PT(613)
     OR ROM32_INSTR_PT(615) OR ROM32_INSTR_PT(621)
     OR ROM32_INSTR_PT(624) OR ROM32_INSTR_PT(626)
     OR ROM32_INSTR_PT(629) OR ROM32_INSTR_PT(630)
     OR ROM32_INSTR_PT(639) OR ROM32_INSTR_PT(640)
     OR ROM32_INSTR_PT(642) OR ROM32_INSTR_PT(643)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(654)
     OR ROM32_INSTR_PT(660) OR ROM32_INSTR_PT(664)
     OR ROM32_INSTR_PT(666) OR ROM32_INSTR_PT(674)
     OR ROM32_INSTR_PT(677) OR ROM32_INSTR_PT(697)
     OR ROM32_INSTR_PT(708) OR ROM32_INSTR_PT(719)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(729)
     OR ROM32_INSTR_PT(731) OR ROM32_INSTR_PT(736)
     OR ROM32_INSTR_PT(751) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(755) OR ROM32_INSTR_PT(762)
     OR ROM32_INSTR_PT(763) OR ROM32_INSTR_PT(770)
     OR ROM32_INSTR_PT(792) OR ROM32_INSTR_PT(805)
     OR ROM32_INSTR_PT(812) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(829) OR ROM32_INSTR_PT(854)
     OR ROM32_INSTR_PT(855) OR ROM32_INSTR_PT(862)
     OR ROM32_INSTR_PT(870) OR ROM32_INSTR_PT(878)
    );
MQQ1884:TEMPLATE(29) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(4)
     OR ROM32_INSTR_PT(5) OR ROM32_INSTR_PT(6)
     OR ROM32_INSTR_PT(7) OR ROM32_INSTR_PT(8)
     OR ROM32_INSTR_PT(9) OR ROM32_INSTR_PT(10)
     OR ROM32_INSTR_PT(13) OR ROM32_INSTR_PT(14)
     OR ROM32_INSTR_PT(16) OR ROM32_INSTR_PT(17)
     OR ROM32_INSTR_PT(23) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(27) OR ROM32_INSTR_PT(30)
     OR ROM32_INSTR_PT(37) OR ROM32_INSTR_PT(41)
     OR ROM32_INSTR_PT(49) OR ROM32_INSTR_PT(51)
     OR ROM32_INSTR_PT(52) OR ROM32_INSTR_PT(53)
     OR ROM32_INSTR_PT(59) OR ROM32_INSTR_PT(63)
     OR ROM32_INSTR_PT(66) OR ROM32_INSTR_PT(67)
     OR ROM32_INSTR_PT(73) OR ROM32_INSTR_PT(74)
     OR ROM32_INSTR_PT(77) OR ROM32_INSTR_PT(78)
     OR ROM32_INSTR_PT(84) OR ROM32_INSTR_PT(87)
     OR ROM32_INSTR_PT(90) OR ROM32_INSTR_PT(93)
     OR ROM32_INSTR_PT(97) OR ROM32_INSTR_PT(99)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(103)
     OR ROM32_INSTR_PT(106) OR ROM32_INSTR_PT(114)
     OR ROM32_INSTR_PT(115) OR ROM32_INSTR_PT(116)
     OR ROM32_INSTR_PT(117) OR ROM32_INSTR_PT(118)
     OR ROM32_INSTR_PT(124) OR ROM32_INSTR_PT(127)
     OR ROM32_INSTR_PT(130) OR ROM32_INSTR_PT(131)
     OR ROM32_INSTR_PT(132) OR ROM32_INSTR_PT(134)
     OR ROM32_INSTR_PT(135) OR ROM32_INSTR_PT(139)
     OR ROM32_INSTR_PT(148) OR ROM32_INSTR_PT(153)
     OR ROM32_INSTR_PT(159) OR ROM32_INSTR_PT(164)
     OR ROM32_INSTR_PT(169) OR ROM32_INSTR_PT(171)
     OR ROM32_INSTR_PT(172) OR ROM32_INSTR_PT(181)
     OR ROM32_INSTR_PT(183) OR ROM32_INSTR_PT(184)
     OR ROM32_INSTR_PT(187) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(200) OR ROM32_INSTR_PT(204)
     OR ROM32_INSTR_PT(205) OR ROM32_INSTR_PT(212)
     OR ROM32_INSTR_PT(216) OR ROM32_INSTR_PT(219)
     OR ROM32_INSTR_PT(220) OR ROM32_INSTR_PT(223)
     OR ROM32_INSTR_PT(227) OR ROM32_INSTR_PT(229)
     OR ROM32_INSTR_PT(232) OR ROM32_INSTR_PT(235)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(241)
     OR ROM32_INSTR_PT(244) OR ROM32_INSTR_PT(250)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(256)
     OR ROM32_INSTR_PT(259) OR ROM32_INSTR_PT(260)
     OR ROM32_INSTR_PT(261) OR ROM32_INSTR_PT(264)
     OR ROM32_INSTR_PT(267) OR ROM32_INSTR_PT(269)
     OR ROM32_INSTR_PT(270) OR ROM32_INSTR_PT(271)
     OR ROM32_INSTR_PT(273) OR ROM32_INSTR_PT(274)
     OR ROM32_INSTR_PT(275) OR ROM32_INSTR_PT(280)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(282)
     OR ROM32_INSTR_PT(284) OR ROM32_INSTR_PT(288)
     OR ROM32_INSTR_PT(289) OR ROM32_INSTR_PT(290)
     OR ROM32_INSTR_PT(293) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(306) OR ROM32_INSTR_PT(309)
     OR ROM32_INSTR_PT(310) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(322)
     OR ROM32_INSTR_PT(323) OR ROM32_INSTR_PT(328)
     OR ROM32_INSTR_PT(337) OR ROM32_INSTR_PT(348)
     OR ROM32_INSTR_PT(361) OR ROM32_INSTR_PT(371)
     OR ROM32_INSTR_PT(374) OR ROM32_INSTR_PT(378)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(383) OR ROM32_INSTR_PT(387)
     OR ROM32_INSTR_PT(390) OR ROM32_INSTR_PT(392)
     OR ROM32_INSTR_PT(393) OR ROM32_INSTR_PT(398)
     OR ROM32_INSTR_PT(400) OR ROM32_INSTR_PT(401)
     OR ROM32_INSTR_PT(406) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(411) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(416)
     OR ROM32_INSTR_PT(419) OR ROM32_INSTR_PT(421)
     OR ROM32_INSTR_PT(425) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(428) OR ROM32_INSTR_PT(433)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(435)
     OR ROM32_INSTR_PT(436) OR ROM32_INSTR_PT(437)
     OR ROM32_INSTR_PT(438) OR ROM32_INSTR_PT(441)
     OR ROM32_INSTR_PT(443) OR ROM32_INSTR_PT(451)
     OR ROM32_INSTR_PT(452) OR ROM32_INSTR_PT(465)
     OR ROM32_INSTR_PT(475) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(481)
     OR ROM32_INSTR_PT(482) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(494) OR ROM32_INSTR_PT(495)
     OR ROM32_INSTR_PT(501) OR ROM32_INSTR_PT(502)
     OR ROM32_INSTR_PT(506) OR ROM32_INSTR_PT(507)
     OR ROM32_INSTR_PT(508) OR ROM32_INSTR_PT(509)
     OR ROM32_INSTR_PT(511) OR ROM32_INSTR_PT(517)
     OR ROM32_INSTR_PT(519) OR ROM32_INSTR_PT(520)
     OR ROM32_INSTR_PT(522) OR ROM32_INSTR_PT(524)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(531)
     OR ROM32_INSTR_PT(532) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(535) OR ROM32_INSTR_PT(543)
     OR ROM32_INSTR_PT(544) OR ROM32_INSTR_PT(547)
     OR ROM32_INSTR_PT(550) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(556)
     OR ROM32_INSTR_PT(557) OR ROM32_INSTR_PT(558)
     OR ROM32_INSTR_PT(562) OR ROM32_INSTR_PT(563)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(568)
     OR ROM32_INSTR_PT(570) OR ROM32_INSTR_PT(574)
     OR ROM32_INSTR_PT(575) OR ROM32_INSTR_PT(578)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(580)
     OR ROM32_INSTR_PT(581) OR ROM32_INSTR_PT(582)
     OR ROM32_INSTR_PT(584) OR ROM32_INSTR_PT(585)
     OR ROM32_INSTR_PT(587) OR ROM32_INSTR_PT(590)
     OR ROM32_INSTR_PT(595) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(601)
     OR ROM32_INSTR_PT(602) OR ROM32_INSTR_PT(609)
     OR ROM32_INSTR_PT(612) OR ROM32_INSTR_PT(622)
     OR ROM32_INSTR_PT(624) OR ROM32_INSTR_PT(625)
     OR ROM32_INSTR_PT(626) OR ROM32_INSTR_PT(629)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(634)
     OR ROM32_INSTR_PT(638) OR ROM32_INSTR_PT(639)
     OR ROM32_INSTR_PT(640) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(664) OR ROM32_INSTR_PT(666)
     OR ROM32_INSTR_PT(677) OR ROM32_INSTR_PT(684)
     OR ROM32_INSTR_PT(693) OR ROM32_INSTR_PT(697)
     OR ROM32_INSTR_PT(719) OR ROM32_INSTR_PT(726)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(736)
     OR ROM32_INSTR_PT(751) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(755) OR ROM32_INSTR_PT(762)
     OR ROM32_INSTR_PT(770) OR ROM32_INSTR_PT(792)
     OR ROM32_INSTR_PT(829) OR ROM32_INSTR_PT(845)
     OR ROM32_INSTR_PT(853) OR ROM32_INSTR_PT(855)
     OR ROM32_INSTR_PT(862) OR ROM32_INSTR_PT(870)
    );
MQQ1885:TEMPLATE(30) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(4)
     OR ROM32_INSTR_PT(6) OR ROM32_INSTR_PT(8)
     OR ROM32_INSTR_PT(9) OR ROM32_INSTR_PT(13)
     OR ROM32_INSTR_PT(16) OR ROM32_INSTR_PT(17)
     OR ROM32_INSTR_PT(20) OR ROM32_INSTR_PT(26)
     OR ROM32_INSTR_PT(32) OR ROM32_INSTR_PT(37)
     OR ROM32_INSTR_PT(41) OR ROM32_INSTR_PT(45)
     OR ROM32_INSTR_PT(49) OR ROM32_INSTR_PT(50)
     OR ROM32_INSTR_PT(51) OR ROM32_INSTR_PT(52)
     OR ROM32_INSTR_PT(55) OR ROM32_INSTR_PT(59)
     OR ROM32_INSTR_PT(63) OR ROM32_INSTR_PT(66)
     OR ROM32_INSTR_PT(67) OR ROM32_INSTR_PT(73)
     OR ROM32_INSTR_PT(74) OR ROM32_INSTR_PT(77)
     OR ROM32_INSTR_PT(78) OR ROM32_INSTR_PT(79)
     OR ROM32_INSTR_PT(80) OR ROM32_INSTR_PT(84)
     OR ROM32_INSTR_PT(85) OR ROM32_INSTR_PT(87)
     OR ROM32_INSTR_PT(90) OR ROM32_INSTR_PT(92)
     OR ROM32_INSTR_PT(99) OR ROM32_INSTR_PT(100)
     OR ROM32_INSTR_PT(103) OR ROM32_INSTR_PT(105)
     OR ROM32_INSTR_PT(106) OR ROM32_INSTR_PT(111)
     OR ROM32_INSTR_PT(114) OR ROM32_INSTR_PT(115)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(117)
     OR ROM32_INSTR_PT(118) OR ROM32_INSTR_PT(119)
     OR ROM32_INSTR_PT(122) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(127) OR ROM32_INSTR_PT(130)
     OR ROM32_INSTR_PT(134) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(139) OR ROM32_INSTR_PT(142)
     OR ROM32_INSTR_PT(148) OR ROM32_INSTR_PT(153)
     OR ROM32_INSTR_PT(169) OR ROM32_INSTR_PT(171)
     OR ROM32_INSTR_PT(176) OR ROM32_INSTR_PT(179)
     OR ROM32_INSTR_PT(180) OR ROM32_INSTR_PT(181)
     OR ROM32_INSTR_PT(183) OR ROM32_INSTR_PT(184)
     OR ROM32_INSTR_PT(186) OR ROM32_INSTR_PT(194)
     OR ROM32_INSTR_PT(200) OR ROM32_INSTR_PT(204)
     OR ROM32_INSTR_PT(209) OR ROM32_INSTR_PT(214)
     OR ROM32_INSTR_PT(215) OR ROM32_INSTR_PT(216)
     OR ROM32_INSTR_PT(219) OR ROM32_INSTR_PT(220)
     OR ROM32_INSTR_PT(222) OR ROM32_INSTR_PT(223)
     OR ROM32_INSTR_PT(224) OR ROM32_INSTR_PT(227)
     OR ROM32_INSTR_PT(229) OR ROM32_INSTR_PT(233)
     OR ROM32_INSTR_PT(238) OR ROM32_INSTR_PT(241)
     OR ROM32_INSTR_PT(250) OR ROM32_INSTR_PT(254)
     OR ROM32_INSTR_PT(256) OR ROM32_INSTR_PT(259)
     OR ROM32_INSTR_PT(260) OR ROM32_INSTR_PT(261)
     OR ROM32_INSTR_PT(264) OR ROM32_INSTR_PT(267)
     OR ROM32_INSTR_PT(269) OR ROM32_INSTR_PT(270)
     OR ROM32_INSTR_PT(272) OR ROM32_INSTR_PT(273)
     OR ROM32_INSTR_PT(274) OR ROM32_INSTR_PT(278)
     OR ROM32_INSTR_PT(280) OR ROM32_INSTR_PT(282)
     OR ROM32_INSTR_PT(283) OR ROM32_INSTR_PT(288)
     OR ROM32_INSTR_PT(293) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(297) OR ROM32_INSTR_PT(299)
     OR ROM32_INSTR_PT(301) OR ROM32_INSTR_PT(303)
     OR ROM32_INSTR_PT(306) OR ROM32_INSTR_PT(313)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(321)
     OR ROM32_INSTR_PT(328) OR ROM32_INSTR_PT(335)
     OR ROM32_INSTR_PT(343) OR ROM32_INSTR_PT(345)
     OR ROM32_INSTR_PT(346) OR ROM32_INSTR_PT(348)
     OR ROM32_INSTR_PT(356) OR ROM32_INSTR_PT(361)
     OR ROM32_INSTR_PT(364) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(368) OR ROM32_INSTR_PT(371)
     OR ROM32_INSTR_PT(373) OR ROM32_INSTR_PT(374)
     OR ROM32_INSTR_PT(379) OR ROM32_INSTR_PT(383)
     OR ROM32_INSTR_PT(390) OR ROM32_INSTR_PT(392)
     OR ROM32_INSTR_PT(393) OR ROM32_INSTR_PT(396)
     OR ROM32_INSTR_PT(400) OR ROM32_INSTR_PT(401)
     OR ROM32_INSTR_PT(406) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(411) OR ROM32_INSTR_PT(412)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(421)
     OR ROM32_INSTR_PT(424) OR ROM32_INSTR_PT(426)
     OR ROM32_INSTR_PT(428) OR ROM32_INSTR_PT(431)
     OR ROM32_INSTR_PT(433) OR ROM32_INSTR_PT(437)
     OR ROM32_INSTR_PT(441) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(459)
     OR ROM32_INSTR_PT(461) OR ROM32_INSTR_PT(475)
     OR ROM32_INSTR_PT(476) OR ROM32_INSTR_PT(478)
     OR ROM32_INSTR_PT(479) OR ROM32_INSTR_PT(481)
     OR ROM32_INSTR_PT(482) OR ROM32_INSTR_PT(490)
     OR ROM32_INSTR_PT(494) OR ROM32_INSTR_PT(495)
     OR ROM32_INSTR_PT(501) OR ROM32_INSTR_PT(502)
     OR ROM32_INSTR_PT(506) OR ROM32_INSTR_PT(507)
     OR ROM32_INSTR_PT(508) OR ROM32_INSTR_PT(509)
     OR ROM32_INSTR_PT(519) OR ROM32_INSTR_PT(520)
     OR ROM32_INSTR_PT(521) OR ROM32_INSTR_PT(522)
     OR ROM32_INSTR_PT(524) OR ROM32_INSTR_PT(534)
     OR ROM32_INSTR_PT(539) OR ROM32_INSTR_PT(544)
     OR ROM32_INSTR_PT(550) OR ROM32_INSTR_PT(552)
     OR ROM32_INSTR_PT(554) OR ROM32_INSTR_PT(555)
     OR ROM32_INSTR_PT(556) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(558) OR ROM32_INSTR_PT(562)
     OR ROM32_INSTR_PT(568) OR ROM32_INSTR_PT(570)
     OR ROM32_INSTR_PT(575) OR ROM32_INSTR_PT(578)
     OR ROM32_INSTR_PT(581) OR ROM32_INSTR_PT(582)
     OR ROM32_INSTR_PT(583) OR ROM32_INSTR_PT(585)
     OR ROM32_INSTR_PT(587) OR ROM32_INSTR_PT(588)
     OR ROM32_INSTR_PT(590) OR ROM32_INSTR_PT(595)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(602)
     OR ROM32_INSTR_PT(603) OR ROM32_INSTR_PT(607)
     OR ROM32_INSTR_PT(609) OR ROM32_INSTR_PT(612)
     OR ROM32_INSTR_PT(615) OR ROM32_INSTR_PT(624)
     OR ROM32_INSTR_PT(626) OR ROM32_INSTR_PT(629)
     OR ROM32_INSTR_PT(630) OR ROM32_INSTR_PT(639)
     OR ROM32_INSTR_PT(640) OR ROM32_INSTR_PT(642)
     OR ROM32_INSTR_PT(644) OR ROM32_INSTR_PT(666)
     OR ROM32_INSTR_PT(677) OR ROM32_INSTR_PT(683)
     OR ROM32_INSTR_PT(685) OR ROM32_INSTR_PT(689)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(711)
     OR ROM32_INSTR_PT(719) OR ROM32_INSTR_PT(720)
     OR ROM32_INSTR_PT(726) OR ROM32_INSTR_PT(728)
     OR ROM32_INSTR_PT(729) OR ROM32_INSTR_PT(736)
     OR ROM32_INSTR_PT(751) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(755) OR ROM32_INSTR_PT(762)
     OR ROM32_INSTR_PT(763) OR ROM32_INSTR_PT(770)
     OR ROM32_INSTR_PT(807) OR ROM32_INSTR_PT(823)
     OR ROM32_INSTR_PT(831) OR ROM32_INSTR_PT(845)
     OR ROM32_INSTR_PT(855) OR ROM32_INSTR_PT(862)
     OR ROM32_INSTR_PT(870));
MQQ1886:TEMPLATE(31) <= 
    (ROM32_INSTR_PT(31) OR ROM32_INSTR_PT(62)
     OR ROM32_INSTR_PT(81) OR ROM32_INSTR_PT(95)
     OR ROM32_INSTR_PT(104) OR ROM32_INSTR_PT(145)
     OR ROM32_INSTR_PT(147) OR ROM32_INSTR_PT(150)
     OR ROM32_INSTR_PT(162) OR ROM32_INSTR_PT(175)
     OR ROM32_INSTR_PT(185) OR ROM32_INSTR_PT(187)
     OR ROM32_INSTR_PT(208) OR ROM32_INSTR_PT(210)
     OR ROM32_INSTR_PT(225) OR ROM32_INSTR_PT(228)
     OR ROM32_INSTR_PT(230) OR ROM32_INSTR_PT(232)
     OR ROM32_INSTR_PT(235) OR ROM32_INSTR_PT(245)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(279)
     OR ROM32_INSTR_PT(285) OR ROM32_INSTR_PT(292)
     OR ROM32_INSTR_PT(302) OR ROM32_INSTR_PT(307)
     OR ROM32_INSTR_PT(312) OR ROM32_INSTR_PT(325)
     OR ROM32_INSTR_PT(329) OR ROM32_INSTR_PT(338)
     OR ROM32_INSTR_PT(378) OR ROM32_INSTR_PT(398)
     OR ROM32_INSTR_PT(416) OR ROM32_INSTR_PT(419)
     OR ROM32_INSTR_PT(463) OR ROM32_INSTR_PT(489)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(629)
     OR ROM32_INSTR_PT(632) OR ROM32_INSTR_PT(640)
     OR ROM32_INSTR_PT(641) OR ROM32_INSTR_PT(653)
     OR ROM32_INSTR_PT(672) OR ROM32_INSTR_PT(720)
     OR ROM32_INSTR_PT(728) OR ROM32_INSTR_PT(751)
     OR ROM32_INSTR_PT(752) OR ROM32_INSTR_PT(753)
     OR ROM32_INSTR_PT(759) OR ROM32_INSTR_PT(774)
     OR ROM32_INSTR_PT(787) OR ROM32_INSTR_PT(803)
     OR ROM32_INSTR_PT(807) OR ROM32_INSTR_PT(823)
    );
MQQ1887:UCODE_END <= 
    (ROM32_INSTR_PT(198) OR ROM32_INSTR_PT(201)
     OR ROM32_INSTR_PT(213) OR ROM32_INSTR_PT(384)
     OR ROM32_INSTR_PT(438) OR ROM32_INSTR_PT(440)
     OR ROM32_INSTR_PT(450) OR ROM32_INSTR_PT(513)
     OR ROM32_INSTR_PT(515) OR ROM32_INSTR_PT(528)
     OR ROM32_INSTR_PT(541) OR ROM32_INSTR_PT(548)
     OR ROM32_INSTR_PT(553) OR ROM32_INSTR_PT(559)
     OR ROM32_INSTR_PT(567) OR ROM32_INSTR_PT(573)
     OR ROM32_INSTR_PT(576) OR ROM32_INSTR_PT(580)
     OR ROM32_INSTR_PT(589) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(600) OR ROM32_INSTR_PT(601)
     OR ROM32_INSTR_PT(619) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(668) OR ROM32_INSTR_PT(674)
     OR ROM32_INSTR_PT(688) OR ROM32_INSTR_PT(694)
     OR ROM32_INSTR_PT(699) OR ROM32_INSTR_PT(702)
     OR ROM32_INSTR_PT(709) OR ROM32_INSTR_PT(714)
     OR ROM32_INSTR_PT(733) OR ROM32_INSTR_PT(778)
     OR ROM32_INSTR_PT(784) OR ROM32_INSTR_PT(812)
     OR ROM32_INSTR_PT(818) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(821) OR ROM32_INSTR_PT(824)
     OR ROM32_INSTR_PT(840) OR ROM32_INSTR_PT(843)
     OR ROM32_INSTR_PT(844) OR ROM32_INSTR_PT(847)
     OR ROM32_INSTR_PT(853) OR ROM32_INSTR_PT(878)
    );
MQQ1888:UCODE_END_EARLY <= 
    (ROM32_INSTR_PT(372) OR ROM32_INSTR_PT(389)
     OR ROM32_INSTR_PT(650) OR ROM32_INSTR_PT(673)
     OR ROM32_INSTR_PT(681) OR ROM32_INSTR_PT(687)
     OR ROM32_INSTR_PT(725) OR ROM32_INSTR_PT(734)
     OR ROM32_INSTR_PT(750) OR ROM32_INSTR_PT(754)
     OR ROM32_INSTR_PT(781) OR ROM32_INSTR_PT(782)
     OR ROM32_INSTR_PT(794) OR ROM32_INSTR_PT(796)
     OR ROM32_INSTR_PT(797) OR ROM32_INSTR_PT(802)
     OR ROM32_INSTR_PT(808) OR ROM32_INSTR_PT(813)
     OR ROM32_INSTR_PT(820) OR ROM32_INSTR_PT(827)
     OR ROM32_INSTR_PT(873));
MQQ1889:LOOP_BEGIN <= 
    (ROM32_INSTR_PT(24) OR ROM32_INSTR_PT(55)
     OR ROM32_INSTR_PT(105) OR ROM32_INSTR_PT(124)
     OR ROM32_INSTR_PT(147) OR ROM32_INSTR_PT(211)
     OR ROM32_INSTR_PT(228) OR ROM32_INSTR_PT(230)
     OR ROM32_INSTR_PT(239) OR ROM32_INSTR_PT(245)
     OR ROM32_INSTR_PT(253) OR ROM32_INSTR_PT(304)
     OR ROM32_INSTR_PT(308) OR ROM32_INSTR_PT(314)
     OR ROM32_INSTR_PT(321) OR ROM32_INSTR_PT(345)
     OR ROM32_INSTR_PT(366) OR ROM32_INSTR_PT(374)
     OR ROM32_INSTR_PT(407) OR ROM32_INSTR_PT(408)
     OR ROM32_INSTR_PT(432) OR ROM32_INSTR_PT(448)
     OR ROM32_INSTR_PT(460) OR ROM32_INSTR_PT(483)
     OR ROM32_INSTR_PT(490) OR ROM32_INSTR_PT(495)
     OR ROM32_INSTR_PT(544) OR ROM32_INSTR_PT(557)
     OR ROM32_INSTR_PT(571) OR ROM32_INSTR_PT(586)
     OR ROM32_INSTR_PT(604));
MQQ1890:LOOP_END <= 
    (ROM32_INSTR_PT(149) OR ROM32_INSTR_PT(156)
     OR ROM32_INSTR_PT(372) OR ROM32_INSTR_PT(466)
     OR ROM32_INSTR_PT(492) OR ROM32_INSTR_PT(500)
     OR ROM32_INSTR_PT(564) OR ROM32_INSTR_PT(637)
     OR ROM32_INSTR_PT(648) OR ROM32_INSTR_PT(655)
     OR ROM32_INSTR_PT(679) OR ROM32_INSTR_PT(696)
     OR ROM32_INSTR_PT(743) OR ROM32_INSTR_PT(769)
     OR ROM32_INSTR_PT(773) OR ROM32_INSTR_PT(783)
     OR ROM32_INSTR_PT(793) OR ROM32_INSTR_PT(802)
     OR ROM32_INSTR_PT(809) OR ROM32_INSTR_PT(810)
     OR ROM32_INSTR_PT(848) OR ROM32_INSTR_PT(861)
     OR ROM32_INSTR_PT(874));
MQQ1891:COUNT_SRC(0) <= 
    (ROM32_INSTR_PT(75) OR ROM32_INSTR_PT(744)
     OR ROM32_INSTR_PT(761) OR ROM32_INSTR_PT(875)
     OR ROM32_INSTR_PT(879) OR ROM32_INSTR_PT(880)
     OR ROM32_INSTR_PT(883) OR ROM32_INSTR_PT(890)
     OR ROM32_INSTR_PT(891) OR ROM32_INSTR_PT(892)
    );
MQQ1892:COUNT_SRC(1) <= 
    (ROM32_INSTR_PT(838) OR ROM32_INSTR_PT(875)
     OR ROM32_INSTR_PT(880) OR ROM32_INSTR_PT(882)
     OR ROM32_INSTR_PT(886) OR ROM32_INSTR_PT(891)
     OR ROM32_INSTR_PT(892));
MQQ1893:COUNT_SRC(2) <= 
    (ROM32_INSTR_PT(695) OR ROM32_INSTR_PT(744)
     OR ROM32_INSTR_PT(761) OR ROM32_INSTR_PT(828)
     OR ROM32_INSTR_PT(838) OR ROM32_INSTR_PT(890)
     OR ROM32_INSTR_PT(891) OR ROM32_INSTR_PT(892)
    );
MQQ1894:EXTRT <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(19)
     OR ROM32_INSTR_PT(21) OR ROM32_INSTR_PT(25)
     OR ROM32_INSTR_PT(40) OR ROM32_INSTR_PT(44)
     OR ROM32_INSTR_PT(47) OR ROM32_INSTR_PT(69)
     OR ROM32_INSTR_PT(72) OR ROM32_INSTR_PT(82)
     OR ROM32_INSTR_PT(91) OR ROM32_INSTR_PT(94)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(108)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(121)
     OR ROM32_INSTR_PT(131) OR ROM32_INSTR_PT(133)
     OR ROM32_INSTR_PT(136) OR ROM32_INSTR_PT(139)
     OR ROM32_INSTR_PT(151) OR ROM32_INSTR_PT(152)
     OR ROM32_INSTR_PT(161) OR ROM32_INSTR_PT(164)
     OR ROM32_INSTR_PT(168) OR ROM32_INSTR_PT(188)
     OR ROM32_INSTR_PT(190) OR ROM32_INSTR_PT(197)
     OR ROM32_INSTR_PT(221) OR ROM32_INSTR_PT(234)
     OR ROM32_INSTR_PT(236) OR ROM32_INSTR_PT(247)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(262)
     OR ROM32_INSTR_PT(265) OR ROM32_INSTR_PT(266)
     OR ROM32_INSTR_PT(277) OR ROM32_INSTR_PT(281)
     OR ROM32_INSTR_PT(284) OR ROM32_INSTR_PT(296)
     OR ROM32_INSTR_PT(300) OR ROM32_INSTR_PT(315)
     OR ROM32_INSTR_PT(316) OR ROM32_INSTR_PT(317)
     OR ROM32_INSTR_PT(327) OR ROM32_INSTR_PT(328)
     OR ROM32_INSTR_PT(333) OR ROM32_INSTR_PT(336)
     OR ROM32_INSTR_PT(349) OR ROM32_INSTR_PT(353)
     OR ROM32_INSTR_PT(354) OR ROM32_INSTR_PT(380)
     OR ROM32_INSTR_PT(381) OR ROM32_INSTR_PT(397)
     OR ROM32_INSTR_PT(410) OR ROM32_INSTR_PT(415)
     OR ROM32_INSTR_PT(420) OR ROM32_INSTR_PT(437)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(457)
     OR ROM32_INSTR_PT(461) OR ROM32_INSTR_PT(483)
     OR ROM32_INSTR_PT(493) OR ROM32_INSTR_PT(525)
     OR ROM32_INSTR_PT(529) OR ROM32_INSTR_PT(533)
     OR ROM32_INSTR_PT(536) OR ROM32_INSTR_PT(587)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(592)
     OR ROM32_INSTR_PT(594) OR ROM32_INSTR_PT(623)
     OR ROM32_INSTR_PT(627) OR ROM32_INSTR_PT(636)
     OR ROM32_INSTR_PT(645) OR ROM32_INSTR_PT(656)
     OR ROM32_INSTR_PT(665) OR ROM32_INSTR_PT(667)
     OR ROM32_INSTR_PT(669) OR ROM32_INSTR_PT(671)
     OR ROM32_INSTR_PT(686) OR ROM32_INSTR_PT(701)
     OR ROM32_INSTR_PT(707) OR ROM32_INSTR_PT(712)
     OR ROM32_INSTR_PT(721) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(723) OR ROM32_INSTR_PT(730)
     OR ROM32_INSTR_PT(735) OR ROM32_INSTR_PT(739)
     OR ROM32_INSTR_PT(742) OR ROM32_INSTR_PT(746)
     OR ROM32_INSTR_PT(756) OR ROM32_INSTR_PT(757)
     OR ROM32_INSTR_PT(758) OR ROM32_INSTR_PT(760)
     OR ROM32_INSTR_PT(764) OR ROM32_INSTR_PT(765)
     OR ROM32_INSTR_PT(766) OR ROM32_INSTR_PT(767)
     OR ROM32_INSTR_PT(768) OR ROM32_INSTR_PT(771)
     OR ROM32_INSTR_PT(772) OR ROM32_INSTR_PT(775)
     OR ROM32_INSTR_PT(776) OR ROM32_INSTR_PT(777)
     OR ROM32_INSTR_PT(788) OR ROM32_INSTR_PT(789)
     OR ROM32_INSTR_PT(791) OR ROM32_INSTR_PT(792)
     OR ROM32_INSTR_PT(798) OR ROM32_INSTR_PT(804)
     OR ROM32_INSTR_PT(806) OR ROM32_INSTR_PT(811)
     OR ROM32_INSTR_PT(816) OR ROM32_INSTR_PT(826)
     OR ROM32_INSTR_PT(833) OR ROM32_INSTR_PT(834)
     OR ROM32_INSTR_PT(835) OR ROM32_INSTR_PT(837)
     OR ROM32_INSTR_PT(841) OR ROM32_INSTR_PT(849)
     OR ROM32_INSTR_PT(856) OR ROM32_INSTR_PT(858)
     OR ROM32_INSTR_PT(859) OR ROM32_INSTR_PT(860)
     OR ROM32_INSTR_PT(862) OR ROM32_INSTR_PT(863)
     OR ROM32_INSTR_PT(864) OR ROM32_INSTR_PT(865)
     OR ROM32_INSTR_PT(866) OR ROM32_INSTR_PT(867)
     OR ROM32_INSTR_PT(870) OR ROM32_INSTR_PT(876)
     OR ROM32_INSTR_PT(884) OR ROM32_INSTR_PT(885)
    );
MQQ1895:EXTS1 <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(19)
     OR ROM32_INSTR_PT(21) OR ROM32_INSTR_PT(28)
     OR ROM32_INSTR_PT(36) OR ROM32_INSTR_PT(47)
     OR ROM32_INSTR_PT(58) OR ROM32_INSTR_PT(82)
     OR ROM32_INSTR_PT(91) OR ROM32_INSTR_PT(100)
     OR ROM32_INSTR_PT(107) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(136) OR ROM32_INSTR_PT(137)
     OR ROM32_INSTR_PT(157) OR ROM32_INSTR_PT(167)
     OR ROM32_INSTR_PT(193) OR ROM32_INSTR_PT(197)
     OR ROM32_INSTR_PT(212) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(231) OR ROM32_INSTR_PT(236)
     OR ROM32_INSTR_PT(263) OR ROM32_INSTR_PT(277)
     OR ROM32_INSTR_PT(286) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(296) OR ROM32_INSTR_PT(298)
     OR ROM32_INSTR_PT(315) OR ROM32_INSTR_PT(316)
     OR ROM32_INSTR_PT(317) OR ROM32_INSTR_PT(324)
     OR ROM32_INSTR_PT(327) OR ROM32_INSTR_PT(328)
     OR ROM32_INSTR_PT(330) OR ROM32_INSTR_PT(336)
     OR ROM32_INSTR_PT(346) OR ROM32_INSTR_PT(369)
     OR ROM32_INSTR_PT(380) OR ROM32_INSTR_PT(397)
     OR ROM32_INSTR_PT(410) OR ROM32_INSTR_PT(414)
     OR ROM32_INSTR_PT(438) OR ROM32_INSTR_PT(447)
     OR ROM32_INSTR_PT(457) OR ROM32_INSTR_PT(462)
     OR ROM32_INSTR_PT(470) OR ROM32_INSTR_PT(488)
     OR ROM32_INSTR_PT(493) OR ROM32_INSTR_PT(495)
     OR ROM32_INSTR_PT(499) OR ROM32_INSTR_PT(526)
     OR ROM32_INSTR_PT(542) OR ROM32_INSTR_PT(589)
     OR ROM32_INSTR_PT(594) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(623) OR ROM32_INSTR_PT(627)
     OR ROM32_INSTR_PT(636) OR ROM32_INSTR_PT(645)
     OR ROM32_INSTR_PT(651) OR ROM32_INSTR_PT(656)
     OR ROM32_INSTR_PT(667) OR ROM32_INSTR_PT(669)
     OR ROM32_INSTR_PT(670) OR ROM32_INSTR_PT(675)
     OR ROM32_INSTR_PT(686) OR ROM32_INSTR_PT(691)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(701)
     OR ROM32_INSTR_PT(706) OR ROM32_INSTR_PT(707)
     OR ROM32_INSTR_PT(710) OR ROM32_INSTR_PT(716)
     OR ROM32_INSTR_PT(721) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(730) OR ROM32_INSTR_PT(733)
     OR ROM32_INSTR_PT(739) OR ROM32_INSTR_PT(741)
     OR ROM32_INSTR_PT(742) OR ROM32_INSTR_PT(746)
     OR ROM32_INSTR_PT(756) OR ROM32_INSTR_PT(757)
     OR ROM32_INSTR_PT(758) OR ROM32_INSTR_PT(760)
     OR ROM32_INSTR_PT(764) OR ROM32_INSTR_PT(765)
     OR ROM32_INSTR_PT(767) OR ROM32_INSTR_PT(768)
     OR ROM32_INSTR_PT(771) OR ROM32_INSTR_PT(775)
     OR ROM32_INSTR_PT(776) OR ROM32_INSTR_PT(777)
     OR ROM32_INSTR_PT(779) OR ROM32_INSTR_PT(788)
     OR ROM32_INSTR_PT(789) OR ROM32_INSTR_PT(791)
     OR ROM32_INSTR_PT(798) OR ROM32_INSTR_PT(801)
     OR ROM32_INSTR_PT(804) OR ROM32_INSTR_PT(806)
     OR ROM32_INSTR_PT(811) OR ROM32_INSTR_PT(812)
     OR ROM32_INSTR_PT(816) OR ROM32_INSTR_PT(824)
     OR ROM32_INSTR_PT(826) OR ROM32_INSTR_PT(830)
     OR ROM32_INSTR_PT(832) OR ROM32_INSTR_PT(833)
     OR ROM32_INSTR_PT(835) OR ROM32_INSTR_PT(837)
     OR ROM32_INSTR_PT(841) OR ROM32_INSTR_PT(842)
     OR ROM32_INSTR_PT(843) OR ROM32_INSTR_PT(846)
     OR ROM32_INSTR_PT(847) OR ROM32_INSTR_PT(849)
     OR ROM32_INSTR_PT(850) OR ROM32_INSTR_PT(852)
     OR ROM32_INSTR_PT(858) OR ROM32_INSTR_PT(859)
     OR ROM32_INSTR_PT(863) OR ROM32_INSTR_PT(865)
     OR ROM32_INSTR_PT(867) OR ROM32_INSTR_PT(868)
     OR ROM32_INSTR_PT(877) OR ROM32_INSTR_PT(878)
     OR ROM32_INSTR_PT(888));
MQQ1896:EXTS2 <= 
    (ROM32_INSTR_PT(21) OR ROM32_INSTR_PT(25)
     OR ROM32_INSTR_PT(36) OR ROM32_INSTR_PT(44)
     OR ROM32_INSTR_PT(47) OR ROM32_INSTR_PT(91)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(136)
     OR ROM32_INSTR_PT(137) OR ROM32_INSTR_PT(139)
     OR ROM32_INSTR_PT(152) OR ROM32_INSTR_PT(167)
     OR ROM32_INSTR_PT(178) OR ROM32_INSTR_PT(188)
     OR ROM32_INSTR_PT(191) OR ROM32_INSTR_PT(212)
     OR ROM32_INSTR_PT(217) OR ROM32_INSTR_PT(236)
     OR ROM32_INSTR_PT(295) OR ROM32_INSTR_PT(317)
     OR ROM32_INSTR_PT(327) OR ROM32_INSTR_PT(328)
     OR ROM32_INSTR_PT(330) OR ROM32_INSTR_PT(333)
     OR ROM32_INSTR_PT(336) OR ROM32_INSTR_PT(341)
     OR ROM32_INSTR_PT(344) OR ROM32_INSTR_PT(346)
     OR ROM32_INSTR_PT(354) OR ROM32_INSTR_PT(356)
     OR ROM32_INSTR_PT(369) OR ROM32_INSTR_PT(375)
     OR ROM32_INSTR_PT(381) OR ROM32_INSTR_PT(393)
     OR ROM32_INSTR_PT(410) OR ROM32_INSTR_PT(415)
     OR ROM32_INSTR_PT(429) OR ROM32_INSTR_PT(437)
     OR ROM32_INSTR_PT(438) OR ROM32_INSTR_PT(447)
     OR ROM32_INSTR_PT(451) OR ROM32_INSTR_PT(457)
     OR ROM32_INSTR_PT(470) OR ROM32_INSTR_PT(493)
     OR ROM32_INSTR_PT(518) OR ROM32_INSTR_PT(526)
     OR ROM32_INSTR_PT(530) OR ROM32_INSTR_PT(579)
     OR ROM32_INSTR_PT(587) OR ROM32_INSTR_PT(594)
     OR ROM32_INSTR_PT(599) OR ROM32_INSTR_PT(624)
     OR ROM32_INSTR_PT(627) OR ROM32_INSTR_PT(628)
     OR ROM32_INSTR_PT(651) OR ROM32_INSTR_PT(656)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(706)
     OR ROM32_INSTR_PT(710) OR ROM32_INSTR_PT(714)
     OR ROM32_INSTR_PT(721) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(723) OR ROM32_INSTR_PT(730)
     OR ROM32_INSTR_PT(735) OR ROM32_INSTR_PT(737)
     OR ROM32_INSTR_PT(739) OR ROM32_INSTR_PT(742)
     OR ROM32_INSTR_PT(746) OR ROM32_INSTR_PT(749)
     OR ROM32_INSTR_PT(756) OR ROM32_INSTR_PT(760)
     OR ROM32_INSTR_PT(764) OR ROM32_INSTR_PT(767)
     OR ROM32_INSTR_PT(770) OR ROM32_INSTR_PT(779)
     OR ROM32_INSTR_PT(789) OR ROM32_INSTR_PT(791)
     OR ROM32_INSTR_PT(812) OR ROM32_INSTR_PT(819)
     OR ROM32_INSTR_PT(822) OR ROM32_INSTR_PT(824)
     OR ROM32_INSTR_PT(835) OR ROM32_INSTR_PT(841)
     OR ROM32_INSTR_PT(842) OR ROM32_INSTR_PT(850)
     OR ROM32_INSTR_PT(853) OR ROM32_INSTR_PT(858)
     OR ROM32_INSTR_PT(863) OR ROM32_INSTR_PT(865)
     OR ROM32_INSTR_PT(867) OR ROM32_INSTR_PT(868)
     OR ROM32_INSTR_PT(876) OR ROM32_INSTR_PT(878)
     OR ROM32_INSTR_PT(885));
MQQ1897:EXTS3 <= 
    (ROM32_INSTR_PT(47) OR ROM32_INSTR_PT(58)
     OR ROM32_INSTR_PT(126) OR ROM32_INSTR_PT(133)
     OR ROM32_INSTR_PT(135) OR ROM32_INSTR_PT(168)
     OR ROM32_INSTR_PT(190) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(263) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(333)
     OR ROM32_INSTR_PT(346) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(397) OR ROM32_INSTR_PT(409)
     OR ROM32_INSTR_PT(467) OR ROM32_INSTR_PT(487)
     OR ROM32_INSTR_PT(526) OR ROM32_INSTR_PT(623)
     OR ROM32_INSTR_PT(692) OR ROM32_INSTR_PT(707)
     OR ROM32_INSTR_PT(710) OR ROM32_INSTR_PT(717)
     OR ROM32_INSTR_PT(730) OR ROM32_INSTR_PT(771)
     OR ROM32_INSTR_PT(792) OR ROM32_INSTR_PT(804)
     OR ROM32_INSTR_PT(826) OR ROM32_INSTR_PT(837)
     OR ROM32_INSTR_PT(866) OR ROM32_INSTR_PT(887)
    );
MQQ1898:SEL0_5 <= 
    (ROM32_INSTR_PT(651) OR ROM32_INSTR_PT(714)
    );
MQQ1899:SEL6_10(0) <= 
    (ROM32_INSTR_PT(40) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(83) OR ROM32_INSTR_PT(94)
     OR ROM32_INSTR_PT(108) OR ROM32_INSTR_PT(201)
     OR ROM32_INSTR_PT(212) OR ROM32_INSTR_PT(266)
     OR ROM32_INSTR_PT(384) OR ROM32_INSTR_PT(438)
     OR ROM32_INSTR_PT(440) OR ROM32_INSTR_PT(450)
     OR ROM32_INSTR_PT(512) OR ROM32_INSTR_PT(518)
     OR ROM32_INSTR_PT(528) OR ROM32_INSTR_PT(529)
     OR ROM32_INSTR_PT(536) OR ROM32_INSTR_PT(541)
     OR ROM32_INSTR_PT(548) OR ROM32_INSTR_PT(559)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(572)
     OR ROM32_INSTR_PT(580) OR ROM32_INSTR_PT(599)
     OR ROM32_INSTR_PT(601) OR ROM32_INSTR_PT(618)
     OR ROM32_INSTR_PT(661) OR ROM32_INSTR_PT(693)
     OR ROM32_INSTR_PT(702) OR ROM32_INSTR_PT(784)
     OR ROM32_INSTR_PT(818) OR ROM32_INSTR_PT(853)
    );
MQQ1900:SEL6_10(1) <= 
    (ROM32_INSTR_PT(1) OR ROM32_INSTR_PT(2)
     OR ROM32_INSTR_PT(40) OR ROM32_INSTR_PT(54)
     OR ROM32_INSTR_PT(71) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(80) OR ROM32_INSTR_PT(83)
     OR ROM32_INSTR_PT(94) OR ROM32_INSTR_PT(108)
     OR ROM32_INSTR_PT(121) OR ROM32_INSTR_PT(178)
     OR ROM32_INSTR_PT(182) OR ROM32_INSTR_PT(262)
     OR ROM32_INSTR_PT(266) OR ROM32_INSTR_PT(284)
     OR ROM32_INSTR_PT(334) OR ROM32_INSTR_PT(344)
     OR ROM32_INSTR_PT(346) OR ROM32_INSTR_PT(347)
     OR ROM32_INSTR_PT(351) OR ROM32_INSTR_PT(356)
     OR ROM32_INSTR_PT(375) OR ROM32_INSTR_PT(403)
     OR ROM32_INSTR_PT(427) OR ROM32_INSTR_PT(432)
     OR ROM32_INSTR_PT(455) OR ROM32_INSTR_PT(461)
     OR ROM32_INSTR_PT(483) OR ROM32_INSTR_PT(485)
     OR ROM32_INSTR_PT(529) OR ROM32_INSTR_PT(530)
     OR ROM32_INSTR_PT(536) OR ROM32_INSTR_PT(539)
     OR ROM32_INSTR_PT(579) OR ROM32_INSTR_PT(592)
     OR ROM32_INSTR_PT(651) OR ROM32_INSTR_PT(658)
     OR ROM32_INSTR_PT(691) OR ROM32_INSTR_PT(692)
     OR ROM32_INSTR_PT(703) OR ROM32_INSTR_PT(710)
     OR ROM32_INSTR_PT(714) OR ROM32_INSTR_PT(716)
     OR ROM32_INSTR_PT(723) OR ROM32_INSTR_PT(724)
     OR ROM32_INSTR_PT(732) OR ROM32_INSTR_PT(856)
     OR ROM32_INSTR_PT(862) OR ROM32_INSTR_PT(870)
    );
MQQ1901:SEL11_15(0) <= 
    (ROM32_INSTR_PT(36) OR ROM32_INSTR_PT(133)
     OR ROM32_INSTR_PT(193) OR ROM32_INSTR_PT(231)
     OR ROM32_INSTR_PT(246) OR ROM32_INSTR_PT(286)
     OR ROM32_INSTR_PT(369) OR ROM32_INSTR_PT(381)
     OR ROM32_INSTR_PT(434) OR ROM32_INSTR_PT(444)
     OR ROM32_INSTR_PT(462) OR ROM32_INSTR_PT(589)
     OR ROM32_INSTR_PT(663) OR ROM32_INSTR_PT(733)
     OR ROM32_INSTR_PT(792) OR ROM32_INSTR_PT(825)
    );
MQQ1902:SEL11_15(1) <= 
    (ROM32_INSTR_PT(22) OR ROM32_INSTR_PT(25)
     OR ROM32_INSTR_PT(36) OR ROM32_INSTR_PT(44)
     OR ROM32_INSTR_PT(48) OR ROM32_INSTR_PT(61)
     OR ROM32_INSTR_PT(64) OR ROM32_INSTR_PT(65)
     OR ROM32_INSTR_PT(69) OR ROM32_INSTR_PT(86)
     OR ROM32_INSTR_PT(95) OR ROM32_INSTR_PT(106)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(129)
     OR ROM32_INSTR_PT(131) OR ROM32_INSTR_PT(139)
     OR ROM32_INSTR_PT(140) OR ROM32_INSTR_PT(151)
     OR ROM32_INSTR_PT(160) OR ROM32_INSTR_PT(164)
     OR ROM32_INSTR_PT(188) OR ROM32_INSTR_PT(190)
     OR ROM32_INSTR_PT(193) OR ROM32_INSTR_PT(201)
     OR ROM32_INSTR_PT(221) OR ROM32_INSTR_PT(231)
     OR ROM32_INSTR_PT(234) OR ROM32_INSTR_PT(247)
     OR ROM32_INSTR_PT(251) OR ROM32_INSTR_PT(265)
     OR ROM32_INSTR_PT(281) OR ROM32_INSTR_PT(286)
     OR ROM32_INSTR_PT(300) OR ROM32_INSTR_PT(351)
     OR ROM32_INSTR_PT(354) OR ROM32_INSTR_PT(369)
     OR ROM32_INSTR_PT(384) OR ROM32_INSTR_PT(393)
     OR ROM32_INSTR_PT(415) OR ROM32_INSTR_PT(420)
     OR ROM32_INSTR_PT(429) OR ROM32_INSTR_PT(434)
     OR ROM32_INSTR_PT(437) OR ROM32_INSTR_PT(440)
     OR ROM32_INSTR_PT(450) OR ROM32_INSTR_PT(451)
     OR ROM32_INSTR_PT(462) OR ROM32_INSTR_PT(518)
     OR ROM32_INSTR_PT(523) OR ROM32_INSTR_PT(528)
     OR ROM32_INSTR_PT(545) OR ROM32_INSTR_PT(548)
     OR ROM32_INSTR_PT(559) OR ROM32_INSTR_PT(572)
     OR ROM32_INSTR_PT(587) OR ROM32_INSTR_PT(589)
     OR ROM32_INSTR_PT(591) OR ROM32_INSTR_PT(601)
     OR ROM32_INSTR_PT(618) OR ROM32_INSTR_PT(624)
     OR ROM32_INSTR_PT(631) OR ROM32_INSTR_PT(663)
     OR ROM32_INSTR_PT(665) OR ROM32_INSTR_PT(693)
     OR ROM32_INSTR_PT(702) OR ROM32_INSTR_PT(713)
     OR ROM32_INSTR_PT(714) OR ROM32_INSTR_PT(727)
     OR ROM32_INSTR_PT(780) OR ROM32_INSTR_PT(784)
     OR ROM32_INSTR_PT(801) OR ROM32_INSTR_PT(812)
     OR ROM32_INSTR_PT(819) OR ROM32_INSTR_PT(824)
     OR ROM32_INSTR_PT(839) OR ROM32_INSTR_PT(843)
     OR ROM32_INSTR_PT(847) OR ROM32_INSTR_PT(878)
    );
MQQ1903:SEL16_20(0) <= 
    (ROM32_INSTR_PT(5) OR ROM32_INSTR_PT(133)
     OR ROM32_INSTR_PT(194) OR ROM32_INSTR_PT(254)
     OR ROM32_INSTR_PT(256) OR ROM32_INSTR_PT(353)
     OR ROM32_INSTR_PT(444) OR ROM32_INSTR_PT(533)
     OR ROM32_INSTR_PT(792) OR ROM32_INSTR_PT(825)
    );
MQQ1904:SEL16_20(1) <= 
    (ROM32_INSTR_PT(3) OR ROM32_INSTR_PT(11)
     OR ROM32_INSTR_PT(15) OR ROM32_INSTR_PT(28)
     OR ROM32_INSTR_PT(40) OR ROM32_INSTR_PT(46)
     OR ROM32_INSTR_PT(48) OR ROM32_INSTR_PT(72)
     OR ROM32_INSTR_PT(76) OR ROM32_INSTR_PT(83)
     OR ROM32_INSTR_PT(88) OR ROM32_INSTR_PT(94)
     OR ROM32_INSTR_PT(100) OR ROM32_INSTR_PT(108)
     OR ROM32_INSTR_PT(126) OR ROM32_INSTR_PT(131)
     OR ROM32_INSTR_PT(133) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(140) OR ROM32_INSTR_PT(161)
     OR ROM32_INSTR_PT(164) OR ROM32_INSTR_PT(201)
     OR ROM32_INSTR_PT(204) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(248) OR ROM32_INSTR_PT(265)
     OR ROM32_INSTR_PT(266) OR ROM32_INSTR_PT(277)
     OR ROM32_INSTR_PT(293) OR ROM32_INSTR_PT(298)
     OR ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(320)
     OR ROM32_INSTR_PT(334) OR ROM32_INSTR_PT(351)
     OR ROM32_INSTR_PT(353) OR ROM32_INSTR_PT(359)
     OR ROM32_INSTR_PT(384) OR ROM32_INSTR_PT(397)
     OR ROM32_INSTR_PT(409) OR ROM32_INSTR_PT(420)
     OR ROM32_INSTR_PT(443) OR ROM32_INSTR_PT(444)
     OR ROM32_INSTR_PT(450) OR ROM32_INSTR_PT(467)
     OR ROM32_INSTR_PT(487) OR ROM32_INSTR_PT(495)
     OR ROM32_INSTR_PT(510) OR ROM32_INSTR_PT(523)
     OR ROM32_INSTR_PT(528) OR ROM32_INSTR_PT(529)
     OR ROM32_INSTR_PT(540) OR ROM32_INSTR_PT(548)
     OR ROM32_INSTR_PT(559) OR ROM32_INSTR_PT(560)
     OR ROM32_INSTR_PT(566) OR ROM32_INSTR_PT(571)
     OR ROM32_INSTR_PT(572) OR ROM32_INSTR_PT(600)
     OR ROM32_INSTR_PT(601) OR ROM32_INSTR_PT(609)
     OR ROM32_INSTR_PT(618) OR ROM32_INSTR_PT(631)
     OR ROM32_INSTR_PT(649) OR ROM32_INSTR_PT(661)
     OR ROM32_INSTR_PT(693) OR ROM32_INSTR_PT(702)
     OR ROM32_INSTR_PT(713) OR ROM32_INSTR_PT(766)
     OR ROM32_INSTR_PT(784) OR ROM32_INSTR_PT(792)
     OR ROM32_INSTR_PT(825) OR ROM32_INSTR_PT(836)
    );
MQQ1905:SEL21_25(0) <= 
    (ROM32_INSTR_PT(197));
MQQ1906:SEL21_25(1) <= 
    (ROM32_INSTR_PT(15) OR ROM32_INSTR_PT(28)
     OR ROM32_INSTR_PT(46) OR ROM32_INSTR_PT(48)
     OR ROM32_INSTR_PT(65) OR ROM32_INSTR_PT(76)
     OR ROM32_INSTR_PT(88) OR ROM32_INSTR_PT(140)
     OR ROM32_INSTR_PT(201) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(265) OR ROM32_INSTR_PT(320)
     OR ROM32_INSTR_PT(351) OR ROM32_INSTR_PT(359)
     OR ROM32_INSTR_PT(384) OR ROM32_INSTR_PT(420)
     OR ROM32_INSTR_PT(450) OR ROM32_INSTR_PT(467)
     OR ROM32_INSTR_PT(512) OR ROM32_INSTR_PT(528)
     OR ROM32_INSTR_PT(540) OR ROM32_INSTR_PT(548)
     OR ROM32_INSTR_PT(559) OR ROM32_INSTR_PT(571)
     OR ROM32_INSTR_PT(572) OR ROM32_INSTR_PT(631)
     OR ROM32_INSTR_PT(651) OR ROM32_INSTR_PT(702)
     OR ROM32_INSTR_PT(714) OR ROM32_INSTR_PT(727)
     OR ROM32_INSTR_PT(784));
MQQ1907:SEL26_30 <= 
    (ROM32_INSTR_PT(15) OR ROM32_INSTR_PT(28)
     OR ROM32_INSTR_PT(46) OR ROM32_INSTR_PT(48)
     OR ROM32_INSTR_PT(65) OR ROM32_INSTR_PT(76)
     OR ROM32_INSTR_PT(88) OR ROM32_INSTR_PT(140)
     OR ROM32_INSTR_PT(201) OR ROM32_INSTR_PT(226)
     OR ROM32_INSTR_PT(265) OR ROM32_INSTR_PT(320)
     OR ROM32_INSTR_PT(351) OR ROM32_INSTR_PT(359)
     OR ROM32_INSTR_PT(384) OR ROM32_INSTR_PT(420)
     OR ROM32_INSTR_PT(450) OR ROM32_INSTR_PT(467)
     OR ROM32_INSTR_PT(512) OR ROM32_INSTR_PT(528)
     OR ROM32_INSTR_PT(540) OR ROM32_INSTR_PT(548)
     OR ROM32_INSTR_PT(559) OR ROM32_INSTR_PT(571)
     OR ROM32_INSTR_PT(572) OR ROM32_INSTR_PT(631)
     OR ROM32_INSTR_PT(651) OR ROM32_INSTR_PT(702)
     OR ROM32_INSTR_PT(714) OR ROM32_INSTR_PT(727)
     OR ROM32_INSTR_PT(784));
MQQ1908:SEL31 <= 
    (ROM32_INSTR_PT(15) OR ROM32_INSTR_PT(28)
     OR ROM32_INSTR_PT(61) OR ROM32_INSTR_PT(65)
     OR ROM32_INSTR_PT(76) OR ROM32_INSTR_PT(88)
     OR ROM32_INSTR_PT(140) OR ROM32_INSTR_PT(201)
     OR ROM32_INSTR_PT(265) OR ROM32_INSTR_PT(320)
     OR ROM32_INSTR_PT(346) OR ROM32_INSTR_PT(351)
     OR ROM32_INSTR_PT(356) OR ROM32_INSTR_PT(359)
     OR ROM32_INSTR_PT(384) OR ROM32_INSTR_PT(420)
     OR ROM32_INSTR_PT(450) OR ROM32_INSTR_PT(467)
     OR ROM32_INSTR_PT(540) OR ROM32_INSTR_PT(541)
     OR ROM32_INSTR_PT(559) OR ROM32_INSTR_PT(560)
     OR ROM32_INSTR_PT(572) OR ROM32_INSTR_PT(631)
     OR ROM32_INSTR_PT(651) OR ROM32_INSTR_PT(692)
     OR ROM32_INSTR_PT(702) OR ROM32_INSTR_PT(710)
     OR ROM32_INSTR_PT(714) OR ROM32_INSTR_PT(784)
     OR ROM32_INSTR_PT(818));
MQQ1909:CR_BF2FXM <= 
    (ROM32_INSTR_PT(713));
MQQ1910:SKIP_COND <= 
    (ROM32_INSTR_PT(21) OR ROM32_INSTR_PT(32)
     OR ROM32_INSTR_PT(82) OR ROM32_INSTR_PT(89)
     OR ROM32_INSTR_PT(91) OR ROM32_INSTR_PT(127)
     OR ROM32_INSTR_PT(217) OR ROM32_INSTR_PT(295)
     OR ROM32_INSTR_PT(327) OR ROM32_INSTR_PT(328)
     OR ROM32_INSTR_PT(341) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(485) OR ROM32_INSTR_PT(662)
     OR ROM32_INSTR_PT(667) OR ROM32_INSTR_PT(676)
     OR ROM32_INSTR_PT(682) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(736) OR ROM32_INSTR_PT(737)
     OR ROM32_INSTR_PT(738) OR ROM32_INSTR_PT(739)
     OR ROM32_INSTR_PT(740) OR ROM32_INSTR_PT(742)
     OR ROM32_INSTR_PT(747) OR ROM32_INSTR_PT(748)
     OR ROM32_INSTR_PT(749) OR ROM32_INSTR_PT(758)
     OR ROM32_INSTR_PT(770) OR ROM32_INSTR_PT(775)
     OR ROM32_INSTR_PT(776) OR ROM32_INSTR_PT(777)
     OR ROM32_INSTR_PT(786) OR ROM32_INSTR_PT(788)
     OR ROM32_INSTR_PT(789) OR ROM32_INSTR_PT(800)
     OR ROM32_INSTR_PT(811) OR ROM32_INSTR_PT(814)
     OR ROM32_INSTR_PT(815) OR ROM32_INSTR_PT(816)
     OR ROM32_INSTR_PT(822) OR ROM32_INSTR_PT(842)
     OR ROM32_INSTR_PT(858) OR ROM32_INSTR_PT(865)
    );
MQQ1911:SKIP_ZERO <= 
    (ROM32_INSTR_PT(318) OR ROM32_INSTR_PT(349)
     OR ROM32_INSTR_PT(432) OR ROM32_INSTR_PT(457)
     OR ROM32_INSTR_PT(483) OR ROM32_INSTR_PT(671)
     OR ROM32_INSTR_PT(712));
MQQ1912:LOOP_ADDR(0) <= 
    (ROM32_INSTR_PT(19) OR ROM32_INSTR_PT(36)
     OR ROM32_INSTR_PT(58) OR ROM32_INSTR_PT(315)
     OR ROM32_INSTR_PT(316) OR ROM32_INSTR_PT(349)
     OR ROM32_INSTR_PT(369) OR ROM32_INSTR_PT(457)
     OR ROM32_INSTR_PT(623) OR ROM32_INSTR_PT(627)
     OR ROM32_INSTR_PT(656) OR ROM32_INSTR_PT(671)
     OR ROM32_INSTR_PT(712) OR ROM32_INSTR_PT(721)
     OR ROM32_INSTR_PT(730) OR ROM32_INSTR_PT(742)
     OR ROM32_INSTR_PT(760) OR ROM32_INSTR_PT(771)
     OR ROM32_INSTR_PT(777) OR ROM32_INSTR_PT(798)
     OR ROM32_INSTR_PT(837) OR ROM32_INSTR_PT(863)
     OR ROM32_INSTR_PT(865));
MQQ1913:LOOP_ADDR(1) <= 
    (ROM32_INSTR_PT(315) OR ROM32_INSTR_PT(525)
     OR ROM32_INSTR_PT(623) OR ROM32_INSTR_PT(627)
     OR ROM32_INSTR_PT(656) OR ROM32_INSTR_PT(712)
     OR ROM32_INSTR_PT(721) OR ROM32_INSTR_PT(730)
     OR ROM32_INSTR_PT(742) OR ROM32_INSTR_PT(777)
     OR ROM32_INSTR_PT(837) OR ROM32_INSTR_PT(858)
     OR ROM32_INSTR_PT(865));
MQQ1914:LOOP_ADDR(2) <= 
    (ROM32_INSTR_PT(58) OR ROM32_INSTR_PT(457)
     OR ROM32_INSTR_PT(717) OR ROM32_INSTR_PT(740)
     OR ROM32_INSTR_PT(747) OR ROM32_INSTR_PT(887)
    );
MQQ1915:LOOP_ADDR(3) <= 
    (ROM32_INSTR_PT(19) OR ROM32_INSTR_PT(58)
     OR ROM32_INSTR_PT(136) OR ROM32_INSTR_PT(316)
     OR ROM32_INSTR_PT(414) OR ROM32_INSTR_PT(457)
     OR ROM32_INSTR_PT(623) OR ROM32_INSTR_PT(706)
     OR ROM32_INSTR_PT(722) OR ROM32_INSTR_PT(730)
     OR ROM32_INSTR_PT(756) OR ROM32_INSTR_PT(760)
     OR ROM32_INSTR_PT(771) OR ROM32_INSTR_PT(798)
     OR ROM32_INSTR_PT(837) OR ROM32_INSTR_PT(864)
     OR ROM32_INSTR_PT(865));
MQQ1916:LOOP_ADDR(4) <= 
    (ROM32_INSTR_PT(19) OR ROM32_INSTR_PT(36)
     OR ROM32_INSTR_PT(58) OR ROM32_INSTR_PT(136)
     OR ROM32_INSTR_PT(315) OR ROM32_INSTR_PT(349)
     OR ROM32_INSTR_PT(369) OR ROM32_INSTR_PT(410)
     OR ROM32_INSTR_PT(457) OR ROM32_INSTR_PT(470)
     OR ROM32_INSTR_PT(717) OR ROM32_INSTR_PT(740)
     OR ROM32_INSTR_PT(742) OR ROM32_INSTR_PT(747)
     OR ROM32_INSTR_PT(777) OR ROM32_INSTR_PT(837)
     OR ROM32_INSTR_PT(863) OR ROM32_INSTR_PT(865)
    );
MQQ1917:LOOP_ADDR(5) <= 
    (ROM32_INSTR_PT(36) OR ROM32_INSTR_PT(58)
     OR ROM32_INSTR_PT(315) OR ROM32_INSTR_PT(623)
     OR ROM32_INSTR_PT(656) OR ROM32_INSTR_PT(671)
     OR ROM32_INSTR_PT(721) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(735) OR ROM32_INSTR_PT(756)
     OR ROM32_INSTR_PT(764) OR ROM32_INSTR_PT(771)
     OR ROM32_INSTR_PT(798) OR ROM32_INSTR_PT(863)
    );
MQQ1918:LOOP_ADDR(6) <= 
    (ROM32_INSTR_PT(36) OR ROM32_INSTR_PT(136)
     OR ROM32_INSTR_PT(315) OR ROM32_INSTR_PT(316)
     OR ROM32_INSTR_PT(369) OR ROM32_INSTR_PT(380)
     OR ROM32_INSTR_PT(457) OR ROM32_INSTR_PT(470)
     OR ROM32_INSTR_PT(623) OR ROM32_INSTR_PT(671)
     OR ROM32_INSTR_PT(721) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(740) OR ROM32_INSTR_PT(742)
     OR ROM32_INSTR_PT(756) OR ROM32_INSTR_PT(760)
     OR ROM32_INSTR_PT(837) OR ROM32_INSTR_PT(858)
     OR ROM32_INSTR_PT(887));
MQQ1919:LOOP_ADDR(7) <= 
    (ROM32_INSTR_PT(19) OR ROM32_INSTR_PT(36)
     OR ROM32_INSTR_PT(58) OR ROM32_INSTR_PT(316)
     OR ROM32_INSTR_PT(349) OR ROM32_INSTR_PT(380)
     OR ROM32_INSTR_PT(410) OR ROM32_INSTR_PT(414)
     OR ROM32_INSTR_PT(623) OR ROM32_INSTR_PT(627)
     OR ROM32_INSTR_PT(721) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(730) OR ROM32_INSTR_PT(740)
     OR ROM32_INSTR_PT(742) OR ROM32_INSTR_PT(765)
     OR ROM32_INSTR_PT(771) OR ROM32_INSTR_PT(826)
     OR ROM32_INSTR_PT(865));
MQQ1920:LOOP_ADDR(8) <= 
    (ROM32_INSTR_PT(136) OR ROM32_INSTR_PT(410)
     OR ROM32_INSTR_PT(414) OR ROM32_INSTR_PT(457)
     OR ROM32_INSTR_PT(470) OR ROM32_INSTR_PT(488)
     OR ROM32_INSTR_PT(706) OR ROM32_INSTR_PT(722)
     OR ROM32_INSTR_PT(730) OR ROM32_INSTR_PT(740)
     OR ROM32_INSTR_PT(742) OR ROM32_INSTR_PT(747)
     OR ROM32_INSTR_PT(756) OR ROM32_INSTR_PT(863)
     OR ROM32_INSTR_PT(887));
MQQ1921:LOOP_ADDR(9) <= 
    (ROM32_INSTR_PT(19) OR ROM32_INSTR_PT(36)
     OR ROM32_INSTR_PT(58) OR ROM32_INSTR_PT(191)
     OR ROM32_INSTR_PT(316) OR ROM32_INSTR_PT(349)
     OR ROM32_INSTR_PT(369) OR ROM32_INSTR_PT(525)
     OR ROM32_INSTR_PT(623) OR ROM32_INSTR_PT(671)
     OR ROM32_INSTR_PT(717) OR ROM32_INSTR_PT(721)
     OR ROM32_INSTR_PT(760) OR ROM32_INSTR_PT(771)
     OR ROM32_INSTR_PT(777) OR ROM32_INSTR_PT(837)
     OR ROM32_INSTR_PT(887));
MQQ1922:LOOP_INIT(0) <= 
    (ROM32_INSTR_PT(168) OR ROM32_INSTR_PT(236)
     OR ROM32_INSTR_PT(315) OR ROM32_INSTR_PT(366)
     OR ROM32_INSTR_PT(397) OR ROM32_INSTR_PT(686)
     OR ROM32_INSTR_PT(717) OR ROM32_INSTR_PT(776)
     OR ROM32_INSTR_PT(788) OR ROM32_INSTR_PT(811)
     OR ROM32_INSTR_PT(816) OR ROM32_INSTR_PT(864)
    );
MQQ1923:LOOP_INIT(1) <= 
    (ROM32_INSTR_PT(893));
MQQ1924:LOOP_INIT(2) <= 
    (ROM32_INSTR_PT(168) OR ROM32_INSTR_PT(776)
     OR ROM32_INSTR_PT(811));
MQQ1925:EP <= 
    (ROM32_INSTR_PT(44) OR ROM32_INSTR_PT(61)
     OR ROM32_INSTR_PT(116) OR ROM32_INSTR_PT(135)
     OR ROM32_INSTR_PT(277) OR ROM32_INSTR_PT(293)
     OR ROM32_INSTR_PT(354) OR ROM32_INSTR_PT(393)
     OR ROM32_INSTR_PT(397) OR ROM32_INSTR_PT(429)
     OR ROM32_INSTR_PT(437) OR ROM32_INSTR_PT(443)
     OR ROM32_INSTR_PT(523) OR ROM32_INSTR_PT(560)
    );

end generate;
rom_addr_d  <=  rom_addr;
rom_data  <=  template & ucode_end & ucode_end_early & loop_begin & loop_end & count_src & extRT & extS1 & extS2 & extS3 &
            sel0_5 & sel6_10 & sel11_15 & sel16_20 & sel21_25 & sel26_30 & sel31 & cr_bf2fxm & skip_cond & skip_zero & loop_addr & loop_init & ep;
rom_addr_latch: tri_rlmreg_p
  generic map (width => rom_addr_l2'length, init => 0, needs_sreset => 0, expand_type => expand_type)
  port map (vd      => vdd,
            gd      => gnd,
            nclk    => nclk,
            act     => rom_act,
            thold_b => pc_iu_func_sl_thold_0_b,
            sg      => pc_iu_sg_0,
            forcee => forcee,
            delay_lclkr => delay_lclkr,
            mpw1_b      => mpw1_b,
            mpw2_b      => mpw2_b,
            d_mode      => d_mode,
            scin    => siv(rom_addr_offset to rom_addr_offset + rom_addr_l2'length-1),
            scout   => sov(rom_addr_offset to rom_addr_offset + rom_addr_l2'length-1),
            din     => rom_addr_d,
            dout    => rom_addr_l2);
siv(0 TO scan_right) <=  sov(1 to scan_right) & scan_in;
scan_out  <=  sov(0);
END IUQ_UC_ROM;

