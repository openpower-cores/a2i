-- © IBM Corp. 2020
-- Licensed under the Apache License, Version 2.0 (the "License"), as modified by
-- the terms below; you may not use the files in this repository except in
-- compliance with the License as modified.
-- You may obtain a copy of the License at http://www.apache.org/licenses/LICENSE-2.0
--
-- Modified Terms:
--
--    1) For the purpose of the patent license granted to you in Section 3 of the
--    License, the "Work" hereby includes implementations of the work of authorship
--    in physical form.
--
--    2) Notwithstanding any terms to the contrary in the License, any licenses
--    necessary for implementation of the Work that are available from OpenPOWER
--    via the Power ISA End User License Agreement (EULA) are explicitly excluded
--    hereunder, and may be obtained from OpenPOWER under the terms and conditions
--    of the EULA.  
--
-- Unless required by applicable law or agreed to in writing, the reference design
-- distributed under the License is distributed on an "AS IS" BASIS, WITHOUT
-- WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. See the License
-- for the specific language governing permissions and limitations under the License.
-- 
-- Additional rights, including the ability to physically implement a softcore that
-- is compliant with the required sections of the Power ISA Specification, are
-- available at no cost under the terms of the OpenPOWER Power ISA EULA, which can be
-- obtained (along with the Power ISA) here: https://openpowerfoundation.org. 


library ieee; use ieee.std_logic_1164.all ; 
library support;
library ibm;
  use ibm.std_ulogic_support.all; 
  use ibm.std_ulogic_function_support.all; 
  use ibm.std_ulogic_ao_support.all; 
  use ibm.std_ulogic_mux_support.all; 
  use support.power_logic_pkg.all;

ENTITY c_prism_csa42 IS
  GENERIC ( btr : string := "CSA42_A2_A12TH" );
  PORT( 
   A       : IN  std_ulogic;
   B       : IN  std_ulogic;
   C       : IN  std_ulogic;
   D       : IN  std_ulogic;
   KI      : IN  std_ulogic;
   KO      : OUT std_ulogic;
   CAR     : OUT std_ulogic;
   SUM     : OUT std_ulogic;
   vd      : inout power_logic;
   gd      : inout power_logic
  );

-- synopsys translate_off


  -- The following will be used by synthesis for unrolling the vector:
   ATTRIBUTE PIN_BIT_INFORMATION of c_prism_csa42 : entity is
     (
       1  => ("   ","A       ","SAME","PIN_BIT_SCALAR"),
       2  => ("   ","B       ","SAME","PIN_BIT_SCALAR"),
       3  => ("   ","C       ","SAME","PIN_BIT_SCALAR"),
       4  => ("   ","D       ","SAME","PIN_BIT_SCALAR"),
       5  => ("   ","KI      ","SAME","PIN_BIT_SCALAR"),
       6  => ("   ","KO      ","SAME","PIN_BIT_SCALAR"),
       7  => ("   ","CAR     ","SAME","PIN_BIT_SCALAR"),
       8  => ("   ","SUM     ","SAME","PIN_BIT_SCALAR"),
       9  => ("   ","VDD     ","SAME","PIN_BIT_SCALAR"),
       10 => ("   ","VSS     ","SAME","PIN_BIT_SCALAR")
       );
-- synopsys translate_on
END                              c_prism_csa42;

ARCHITECTURE c_prism_csa42 OF c_prism_csa42 IS

 signal s1 : std_ulogic;

BEGIN

  s1    <= b  XOR c  XOR d ;
  sum   <= s1 XOR a  XOR ki;

  car   <= (s1 AND a ) OR
           (s1 AND ki) OR
           (a  AND ki);

  ko   <= (b  AND c ) OR
          (b  AND d ) OR
          (c  AND d );


END;
